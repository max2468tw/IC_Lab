`define CYCLE_TIME 6.0
`ifdef RTL
	`timescale 1ns/1ps
	`include "SA.v"  
`endif
`ifdef GATE
	`timescale 1ns/1ps
	`include "SA_SYN.v"
`endif
module PATTERN(
////output Port
	clk,
	rst_n,
	in_valid,
	in,
////input Port
	out_valid,
	out
);
//Port Declaration
input				out_valid;
input		[3:0]	out;
output reg 			clk;
output reg     		rst_n; 
output reg     		in_valid;
output reg	[3:0] 	in; 
`protected
A8EE9SQ:5DT^<T?YQH^=aO62`:]D=DH2n;E:IkK_McYfR38<^ffeCZJ9I_mp:c?j
TV:5ZG^R[L0jZM6ep_\4FaoGDY6I^?A8>e34jOEf0n@9:Z:ag69b=n2@G@1D2KL>
WHojYG0pT5`SZmpFfIDXf>_n:K1@h_0fX>`lfQ91MUiIZJl>?qRViPUO;][eNa7I
nC`@66F_4:oe6;>j_:VP^=6;R`pA?kDBBhje0PkYghqMSY_W`f7<b[GNho5q\RgU
W=9BcOmmi]XJXm;f^P2]AHDhaMKXFR>14m2J?XSVd[G=\Nm=>l18=NL<YJdh75YZ
4CqDG5C0\Z2XG@AHH_bLhPHRhBI[:QmY<IAWH@_GS6PZ>JX7Cq_O1WMD`M454ZAE
S:77OlV=CCZ:\@iLTU;QPedocHE4Z;09^ap8^?^M;5N:ESHPg?CS[=_ZVCK9S;^q
07MB;WQAAWk@gl;k7NP6IcYVTQ=L2fUhQUchj>L]Ldq<\^nN]fTnSa1og=22:NDk
N1VpbKOcc6o?>XLYXVVRi6[341]d`[3flBcPgEUfPbI\p1Qie2Sl7I_NgX_C>]T`
bHHP0OlQ[jSFOa:c>?;Ya5IBqnR9bn]W3^1eQgBC8WbmA:EZ2V^@NGaaX7@Vj\Iq
1fTibY\_lhdSY>F9EY9lLgIgg>j7cf7gGHXFZ7G]o]@^i698CZi>[kPll[pAO3oe
>aAOLjHBgP0HBK4L7]XLLe6ho3QjbGp=AA19leNon@Z@ZXN1\8BhdI0i9Ye0_`kL
mFI`:AP>ljLJKpF3HU0DlZlH`;;V\E:CmGIDpEM]545H1qW_aPRgZ;XE5;FSYn]e
mf4fPaPlPT]So6XKZ8U=[MEh`9cWoJhi7`:76KJmo\=>QZj<3DCKSq3F6?Q]A?ER
bc8D\ODOF?U2hq]4[ER\dCmO;d]c0o9@2dT776gbG6^4<dNdGfJ>CMV]mUkLbD`Z
;J@?6ORAC:=LAqA9_i3gEX3T=[EPYZ7NkC\nWYUP<WU=kpEJOJmjcBNF[]E2bBB:
XGDOHqZl=gLefjO]7ThDTQfAVp75HmV2Q[kCP@nCRCcBp6FQj1K:YHX;5QW[R43J
ZofL0MLWa4iXeQIgEqXBO>188?:48f]0WMJP^FZhSQh^nkBJkaF=pG^`_S[m9P87
490F_GAc=1\jWo;=kp_OO?YfTTE^mgQW45_DNF?Ja\aB583A5M;^bDQ[M1K1e9Wc
M_OO2V\T=qH2O9b[H<aCHG=0Eg;g\dq;Fe??7pk5hk\:q5hZ9DkkLM[\C<?K[Cb7
T7<RmQD>aj=BFO9PLBWmQqLDaCVQjpaN7?ncL5H5<E7Xc:IK;AFSI::kB@dSSH7\
H3]goG=A]48BCbB^^^kIQE^`X6@T`qg=;2ZP[kn`ZhK82LRNJj@\MooU:;UXWPn;
O6?O0QOdn4=0^7HE[j3H^[H2gnqX\1B>IAp8_I\^[pVATY0G0_0g<AG1aB5:D<a0
_?OF[5OPmHcAJZIRDdhi0cJ@F>Ej?SJYjj@l4CdeOEJ^DWlFW5f]0DdVL>KSMLnS
9h1l`G@Gh5\]A<1U?D4Ro<ImcoSd\c_617@BY?oI>eNC@kjL0VUZ;WK<i]d0BX<^
niReK\baS7H\fi<X@XaEO?PBFK[B?725<4pdJZS`lB5G:961@e9KK9FJdIAfJlRb
?_1f5m<=\^OK[_<F<AO\AaYd8DHW9@iEZJGk<SenoQg=3H2nNMh^\F9cXlNQ`l8@
aVZ9i4;A2VF>kJIDR]NlVj?He9?2kmS:HS3>iJn_B6M=`4?IFdL21l82fF1]I1^L
HVDDVXSlVlBVh2e25[O]jaG2FWHpWI\UWVWR<;W7ZZQ3DfWMAo6D:=U\<bCd[B?>
XP=_ZBEBUXKRa<5bIn\:>J`keWJW_1b=DCS>Ea?bkK\U:Hcn;3InJ1GS>oJ^cMhV
<G6D]RX?]Y<DFg=\@^E`4<0S3KKdK<SjP=KQDJE;1LlZGWUGf`k4YQnbNH=L1WIl
0kQ_K5^KG70fo359Vk[Sp7U50?ODi6EOGia4g9;`FACP7Vn3_NibS:MUAY[_3g2m
SImEkl7::qSR<eSNLiKVQ<``n20gY0bkm5Ha5`?F8`4LiDcff_mVNeX:SQHRKhfd
5;:b`[6R4:[ea4P7Ymi1\lAKaHAlI`2DgHAD[bAJo<J:TU:TXASiXfOXeMQc@UJP
Hn_I2ilIPhQCZXbHTjP2U@V[K]7AR1]B?I[IjZcfO2[RFVN\J^7gM5D?bO^YK:<=
C2qL;6`bVB5D[PAm=NPT9og>RjO_HTK\0>FcCW?a:NTEeZ3OcbRZ6JU48@_b3=Oj
LbHRGB?>giHg<X@9BBaV>5^Q[\Kmii8W1<FJ1HHIoI1?=jM??Vi@?1nnA<J]aCcZ
>2@>lCLmZWkFT;h74Z@eFL529DfnoLZTn>L0A6NDH1^:Tn;Xoae?PJmB^`Wp^H`D
0f_W?[`2;N7`Ng8kF:S72BRcb3:JRdZ0_UNTEgIJ4nI;EXgQ1XGC=O]=f9ehhQ8\
5o]=EI7;:j2:K?1le<N3P?5f^JW;EF]Q1G0>g@7bF:kQ>\MPiRdnbcYma<\ZBMND
2?`hh4lKaLeam2kEkcJ[NM;J;mg\7LW5bU8HSA43GajcP6gQG<<>qe1`7XO8LZ8I
\AnIBMn>M<:U@>nJOkFAR7G4O?\adP[PNheo0AKmBYj;U`L:RM1^S2ah9gY`LPmb
al9<Vg<7Vah;_S84LUjd0d:@C4\Pe`OlRoVG]4`fJnW]0AbOoEcE][47e;c9dhHl
[JfYNoBK:M6OS==cVM9Yl0PJH>LZ;<am2^`^;USm?Jf_opj5cG92N5DR;JNURZk3
K:93M_M^G4Cf`YQ[M<dfAiTJjAcmgAPKnf190b2M3FCRHccI;NjdgX_J4HLo^OI>
BncK6\Tc>aQ31>g<XhgYI;d[D[hcmMSZQlm3[05odG=7V_OEbB:8O8RD<90@V@92
YnT6j6PKR?:B@iRc^?Jj76HVMNV:OQRDn^MM<ep@R0VKGQdb9X4mYc^?W\RoSMWU
=RO_`j8G=OkYd\jWnba1_k90gon>>HG=nfE\7NQk9DHddahfIfWS]nmGSfCGBGU2
M0PeoYlfjlRR;lL4GlkDWmGEQRU[HYT4DHaL@T_>Ma8\1[CHHYloC9TiL>CXiinA
LEIXQgeCT4P2U:cC3@9L65haOoPQEdnp>BLo1i^T;kbe\V3S9_8=o5?TiS<;;=jG
?KE_7HWNbVMF@D7JUcm^BKQ:<8GGKGH45_P>boP:>fFf1V^FfekZ;@Fm6FChhKFo
N`AHmfknEZ@\7BFHImkPV^T=7YN;<b@oUcE]\mBIJa^WiS`inT6Ce?S^;9oD=On;
K;KdZ0JEDl0DJC]3V;mnZY2=qXf]8\b@m>TQibneY=68_N2g[lBP`YQ=9dYWX6mP
;`o7DQiYPCKJo_FHY@oNF2o\\a=5WoOb7blh2YVONMioZZ6BMOoBTKX0Ci4>?MZm
`\j@`7[O>CeEa`C^Y[<NmGU=:BSYeUlBX00aQDkZ5[k79cI=JWN=HdYVOFa[o]jH
iMFgB0UlU<kJ_f2;_qL<hd`T>Jn]JnAKhSf:D^_XVXRHhfia:9HFGlU0UjO0\Z9A
@[L_WMJIn>aP4]G8E:Lb72PU;>V4N9YRCoMkRR0VGmhNRA59hoKRYIZQ1NoRaX0g
9gmCVI8WoPWJTF6\oj7<O]VaTVJa0NWILlna0gGh9icMeT=O8n8TZ[5[Vf]3<S7j
gk9VWnGKiIq;dX4K9`>1b;0_a<U]WlQZL\4\LYbK4cC3gK8]:n<Hhiq=]KO?a15Y
N:j>3[Zeb9V7UEQAT3l=3FJiP5Q8>M7?>RSG=h:0G[Q6bY00C[>h[Uc@:9gFH>A6
m]PSR;KgXBX_B6>=maSX5=I4g4F<_L^6<:JE6YXST[F[RQJnD\nK2Y]ILJZQT@8[
_D_V2e125>kWm2P8XUR?VWP<TGfl:PB2U<GEkeN`>[_6AEMq\O_chj1hPZ<G@n9Q
N=mndS=7k:`CnkCDGoEXdlf2BDKWEAdJ?hg_n\ch;k:?SYKQf\5OSWI5BbUO?]RY
?JWAel>YYkh]^Q0AldKeMHT2LKMBl3^??WmlQdGokI:2^LV^ffABZPlUbcGhe?Mn
X<l\Kk1X\WoV`d\JNR80XfU;PZ[YkKGR_:ghN9Qoq3Mc2gDPDIeHYfS<=<9@g;SV
oHS55DYZ5Z`c@<BgL1DooUlS?oE<V>FQd9j?=T4_8k3O=clO:=\h;@b;U0nf33OH
oW6cOPdL8[S710QkadQ?jn7NM[j4@59i?cb8;;4QYHT[iMFBBEOR\]F\OURm^aT[
9HN9m]=JYgaZb`VhHD8XQR;<L7h<FKi<NqOWecYS3H0b^l4:9<cLSZLd8F<DBhGI
]Ni<5Ca<9]4l6l99^_=gUFJ`Y:AeDe1Vclj85O1`WWT:gV01OJ27c8RkjN3hM;V\
\NccE<]5?B:C]nXjlEUC>WLBdB;S@=njkSehZ\eB<?Vjm9UGGX0<WX7m9U\O5@Y]
Cc9AOnjKOAi4eEU<]P=3U[I\JNq7dg?2KG8HCUCS39?TL7E2_8P2>[_F_UmW^`8d
:Cnf?A:hFCa2Kb^0QUC0mWTY<=;lL=YBnd]PTRSP[5KP1Mo?j[2gMjnBD]T?kSV\
AJQ<L]l:iKY>7gmo7:\T`MEgKc:i@\AQdg32Dd05YN59j@D8=fQYEFFC8j8oB:;G
2d2Kj]^JIQk3AbgnjWopi0QY<WJT[;kfR@U@n2<`\S_MlBOe6GO>TTj]n\Eh8\d_
M[P[0\:gboj]L`hT7kT7EG_O]3L0Pjg59TW<Y:;AZXT9JMk<ijXIcNB>`[<K6;NI
em\4XQ0h1fJd6=>W\MhGIe[C<B9_V]<GLARa3P5`EBV1joM\Wc8[aI<\mj9b\o^n
2GCDWX:lFdC5qCHSN@d]=3Yo44Yh2>do[dU2g86>99II>[H;VBSNY2faC=N;cc`=
]o8IP`ff57d><a^hfA2Jo\H4;\:7ZW?Z@FKmiV5NTNEHF[0PoDBI^EnF[anmlQa^
SGDAj0Od]=LOdIj2YM5AJOaWNENLj=C?n7B>Sa\GLK;80f?46I>B>N[W_6aQPLj=
O3`I`pNDh3jo:Sj`;De8_?jb731VaY;Z<[\=GpGGJJVBg_a>=UjN9a<4nVC_kV=]
Hh>Gnojd5P0hjkWeSDdBP>K;ETfU5hX=cj=dPIobVNm`4S3_MIDCYa:KkY1RFC6f
\caD40eVbWLW9ONS8UJW;IYab;a@@Uc?Nc@O57OGBBmo7K7KC1QN3di`;U^Ub>S0
2lHEYN87a8hK>gg\TOm=ZF2PEoI97hpfP_0VJ4Y:4FM64Z<?@7TbkDQXJNfZ^QU8
Um90^G2N=aaOZ9jZFan8`NZ\R2jfE`\HGJFXY125bcXYBAOUHkQGVCnZfoXbQfm<
VFD`@7c9gc:Y:B]4`>mY_5KdkcHAhBMWJ\9=k`D9`Q[_DQj;VX<]3HF_OQoFHO_f
XBPH?fK;]26g8mEO]a=_CIWqmAUGX<geZS5XM?_7LMbI\9YS=Cl\o4i2JG]PNg_V
GZZV_;Z3Dj9MW8g;]0amn4hb\OO>5fEJc^VKiM[TIe0I>cQ=<5<^08jjMo=6X=9i
1PlFVUQUJLDJf?Kd1\TbIC5R@2I3:gbeFRYSRBYIVVHK@GR06Yao9MfI1@2UgJG9
6V9?RK3go^9_kLYYqmm0kKKG`M<j^V4E7nmoUBJLn0NZPcT]20:=10DN2ZRLclf;
ik^D15o14@_Dnia;5`gOL9:QdI8V06DbLF1eM]<[c;RJ7FgC>=EaSZWHLH`7hI?a
ejIARPCb81@g>nFVKlhjEYH;nPnB:lTYiPIaZ:8_33QH@[3::K4hIYH<`i2_AZ2>
YcLDLMo\0q6JLM>KX7Z2nFfhKH@GI9PY4]iobeUc]f=Q1F`>70oEckCO>:c_bPFl
X5NDj@12;LXUM9\eS8AnXXhERX0bUj74ae<Hl2PQB7@8>HRNLBaQF7hN1T1LUdok
j^\iUcjlDY>TWE;[;H\?KUnA\:U_SdUOhVZOHkmS;1RdL[^JIaaBFgUabDiEbYa=
<CqI?ik8FaceWYm4XGoCBjV>6IjSmZ;cj:ML>PVJil15hnP`F`8Jl1@j^ICgc:Tl
]lZKhZ\mWpS[J4:DpH_\]d`PR@Vag=8;e_>=Hjl?YlK]SQEJqX?YA4Gg9G_?mkJ5
jRFeLma`k]agkW0T_SAichco`a5q1g]HgPapPBWY?9S:>LT>aj@l6eIl6FNab=ip
HbGdZUe`?3Oi>I[5Mcj8EIUMSEapVOc5kA<pf_A0I8NL_iahKEj[oICGWP4GVO75
1g3Yfbi9?UYQp3bn6LBqI<ZT2Kj\@hBA[N:0dL0Wgc8K6k:Q;Xmb3H:?]X8pU\Zb
3\B<6]dWH8:A[YkHG2;DHkB2m1JR:3lBRCkYGkK`ajaJM5LCq[\aVl8?W=Uf??<K
`1d:KdgEf0CH_RY2F=fEiXefa?AmK]g:VKcp;^G:KXEWLjHghhQ;IO;XmYXIRA2c
@bbFQc?nPi^mQQ?G;TYqH0TV:2X3d\J82h;9ebljCOb9^_ikW8m97]0oHOe\:PIF
qd@NTb`S^L^WR@;OSSHgigo3bgbkVLiNMh=qGLPhlB5XMNlgoV_THnM=aESb:VlD
Uh4n66<oo2q3CedZ=qndi:LTd0;3<[dhnki4>[_Eb7d`2>e5YK4DGLo\HU5AKpEk
ko`GQ=VFS^H<mk\5lKUIINHRR`oHT]qe9XNXHjAcB0WONJL7I=RC9TO8KaN6W;gJ
6MpY:MenKeoM[hWUN5[Y3RQlWm?ghHMP`AiB6Em1ZS3BB6@WOp3fC4K>P@^dn?id
5bU>a[BKPRUY3ICYoRY8Qko=5D>ef8h:qGMgNMjZ`ZcGk<=>8jdVAX:FM7ZbC5mf
[fTiV]k4?PonTiWq1n_Y7VhKOSHTFi=OFRBh_KN;UCX`KTlOLT1JJ@[:Qm?K3[qT
^mQU?i<aa>m=WT`Bn1TnAkj4km1J7Do7b`7OPAnV;33W?p:CFkDKqBn2g8QbmTLG
\BiKkaUG:mm@nR53@RoCN`<FQ9kZ2\]WX8B<OV4B[ZA;mL@0BqOBcgk2qCNlK;8Q
W32BZM^7Id`fJG=R]R1D22@_e6WhnXaTgONMHanYVj3F9B:\ULZn<j]X29oCqO_9
gJbpN]gUD6q?a`<`K=]]9RGdPnSFYqUZKUoVni^W5`AeE5oVQVMd4q<ndBCbU?4>
<DK1eX:Jfgh`2clKbZm8?ZbKc^qbaKL\7Tq>GOCSdF8^laL];<TghN8052cckd]F
12BMkAaIkUBefoP50mW5N2:^V_:X;bLpXiZ9B=NODHfXhB4c>KpT\1KR2I_K^cJb
EgN^7YK1SUSPal=@X7:U`7qXe^RDoq2TJ?Lo3U?1g7g4[TdMLdhC3idfj5pcJ6IN
OLp:[aMSgpIQX1d0mnUllZI4?M?76;\bbI<6P<@QnWkL1O5<l2If7Y@2BZEB5?QL
n[HQem159FN7g:10mWUllZI4?M?76;\bbI<6P<@QnWTM3i23YLMYmm6\<3SEUq73
110hl:M:;nndVgQ[ni0oJgG9Bn1^MeC;CoUB>M=I9LEYUQ\m?M<2FZi@c1NeTeaW
4QWl<qJ\:Yb5Mb?\fM3kO>KAUWBLkEo4UM=RYbHcPEg5i5j7MD:UO:e\:13_a;<\
T\YU]5J?@Vi5MT?\fM3kO>KAUWBLkEo4UM=RYbVCP]<B]8Z=>CTAAUi\Gq>WB`ZO
cQ>bL43g@5F>E1?=hEkB<_I2=TBabfVNj[]1`5X7Y<bnYPa0:]JAe@OCO]>JEBR]
TJ=0LKb1HBX>EA?VlC=HkDIO7d:G?AQ\DlSOm;0RcARU8EpF:Lm_^Z023:Alnk7G
Fi3>Q`>X7@L`MCX=\liJDb]`ciM<C\>L^C0FY>AEh=KZh:3D>SNL^ZF23:Alnk7G
Fi3>Q`>X7@L`MCX8BS?XNHTg`B25QeF9ZQq``QVAlh_7_Vo[7TMGSCgLOQ\D2dqK
gM7H`D`TT0iF5hOT`>`f>NQCHdL\YFXqZTgU>?EhHDE=:5BYpX@EneKdp>IZ]U\1
pbLP\k9pMeTXgY2>@?_V5KFc72Ji5iLKdYqL1K1DF38GB6O1S]\U:5APM?gNHHDh
Q@j6_:eCYHN=RPPhk3WbllAp`=NHg5q_aX8?IZG\^Sg8Hcq0:HV3E5Vn2QX_CP26
EI^plJkLYJBabCLQ3b=cX7^S;dlRghVRC1o>7V:Oh;J2Ke1@okEbVc7;SRq;PKC0
63p2Zo^7A[7<RV_GCjNe?OJPCdF\C]JbJ`S`D0A46XnOGfp@?i@HfZ[EN@`efWZC
:]H?ElVV8Tq;P4bBM0\e?4Z5DWi7oGXIZk\8?M4:Rk>bXCpAn5_2dW;9XMDU830Y
Bp8N8L5]9YElATImF3TG0MhZW0og0f:=fgU3q322F47kpC@8U>OA3SUmc@YRjA[l
ec5IHARmK4KLj5DpP^kII8@9oE>JgRi65Q`q=b611hVd>6=b^\TamV5p3]=Ya8hV
eSkCA<pJ4E]ZLfp6QoZB4_==d\>Kh4RTbRZj83:4NaUjY>Q89qM>WODXSl0bT[`i
E`9C<1S<H^;jMbB=;Q@[pCXSESfo::VUYV]HeN<YQiCpR_A?U9p\FTPLBqfmC]f7
E]1ihmo@d;0;fB0a\5p<lIZ=[DW2SKF:fJlaKK;7ngHQ:heL6]S]m4]mOkc`C@SS
9]dd9HH@ffK>jT<2m@q4:DhbD=p]o6Q1Jc9O<noSeeb?jW@\8G0E;[_k5EGA6W:S
IQ2qL;UYG::q1\WQ^k7?7YPM2KBhTj@I3NI`S;OLHIGYKY\0YGp62kkCkN4jW2UM
Shf@SOeP<JUa`@?TX=3dfi4XAgn7k4ffZn92aqMZei47lHQGdE\R`VcP9^q[ZRE6
k9pX2D1CIq1RXdojpZn<GhbcC][]E1K5=jiP<]ka8Y@]m7^KLR@T_@a[mGO[m=U4
LPVUUpj<[W`Yp6E^ZODH=V1DMgmPOg2obCdhq\HK3C^=qhjbF:Eq^UK3L7F3cj\i
BUYIFUn<:OJLTMC8<inGL5<CF3Y7n6GMnMT<;JG=R7bHFJC84DQeKBSdR7F3cj\i
BUYIFUn<:OJLTMC8<inGRgBWMgJ6g0<GBJ>CC8hpLGO`bY:[IYB<dl7CO;R<;^Sm
im\oD3L_K2\JMFm>@X>QCT1<:2`J?cN1WiDI`j9hLTJAmY:@IYB<dl7CO;R<;^Sm
im\oD3L_54\lKPLP;W[d6Yl8mAcq\khjP`lo;eUGYfQH0=7HV]XO03iC[6NkjDA8
BSXO[>BRf<gf:U^4Ee5<R;C8;6Ad\aggW7]:aeUBYfQH0=3Y]]MOSS<R][m_FDR8
W[pT@Q_7@<fnC6@CVLmIl7NXmGNheUIO2V^:e^Z[b7IU55`3fEWRJ:H?IjAZ`Ti9
RfL14LKH7@pZi:cbaLFV0a]=4M^6E`?PeHVBN:>h[jE6fQ\60nFo\`bCmbHEd2CD
GAPF75CTH[mZYJM5:J2\bWc=4M^6E`?PeHVBN:>f>C5jb193Yi5lHTW^A3Z`Pbqe
lY<lXCPSYfG[YEIbhQkVI[I]G;`D=IAN]jQZC<JI27B9?WkOeaZ@K7E\FI1Xa;a6
NB4jXCPSYfG[YEIbhQkVI[I]G;`D=IAKGNUAHG4d2M:n_k]Ke=pf[mC>^k;_aod8
\:Mg^49O91^Anbqb:b:f1PVYA5g_]@1;9\]IeFZ>Safan4MS5qiP>[:YPjjBL4Gm
WaqJ;H<IMFH_4BmQO1ce9oIq>X0f8ibqQa7B3?\qfW__:RpdDE0_Np6J0bW090W\
Y;Rgh\HgpCOi_=>HmE_RalmHOW>NcKk[qo^[D[4Npk]RQB@fboeja9D`Q;4WScJ^
OqPkc>3W0o^=BY4_F`54l8B9ClCD:a1\[c<bSGdSM^=Xn^EJ8@E9SIQ@65NdA[ii
Tl]4Xh4SVY>F9NpHThII6VQ_b0D`[<\=nJYjlH9ZJW\lbG?><CV=gR34PPdo``Ed
kIo97@[>4RJ<2KYKVPgI[OO40l=ChCm=1gKq0aGVH6HRZX\39j3SoCk8nRm_eBo^
6Of0OI9KhhaWNeDDeDoFGe2F\YHTRCaH?o83e:J<PFEV:dC`4CDHQEd1BT`;q3Mc
2mBFjTcQoUZUFd37RfaO:=\kDS`_oINbQ_i[E[f:oWB:dXAk5D_j<iCg^OJdV?]G
OQA5lE5Xg0i0bVOUP`mD__9p__iieh>B\4C4B9cXhj6oeO2?T0kcAF6A86H>CiV2
S[U^A;W?IeO_oSjH>IMgH@O45dJa[`R0]0i6<74d:7=KpldRW=@8V?O2SPKJCh4f
ejnL^ZfM0h1:6];lLoE]lY3NjDV:j=JGbfGYc=;EVkAj1KHQa[l8UbP7C@Wb73<:
p=9;:L];JZKjEg1J6@KlGL7?B\72g:I251]C?b6e>^`F_FN>P9?lLHDXCcIMM?1l
L3=KYGAICWEm;?c0HK;T7qg5PFc;Z6?gOBE52J9kfU>e\>CkYk_d^5b2>DPnnnHA
W>V0hApGd^mB@k>eE:Mf9N?oDIfPKcGkDH4]Wi5oo;_7D9CZ<6`7LCfdVF3Ik0RY
3@KJ_d]965TP8=TnZZeOC@2hckjPdM\p]UC]fdj=`m1H3NLMNdmS1V;DZi^LJfI7
7d@iRWGeaT<kLhLKoP:HHH:]EoQTU49>MN:o>1XXdM8UhH>EE0HFY1pSIGB:=<8n
fcI9E5WJlMK1K?U3j62_66Ln<Z[7Rh:=Nm?e54@8Gj>^[[6L06IAGiAnOic[2]F=
TJQd`TJp_aDTAAogaHOnlUU1P@Wn>F[`51d\coHh8mZhT>OL<l7k4G6Dj20?\DVV
VL>FJ3oeMfAAn0?MiEK:q1YIZ`dImLJW2Ha=nEUG2UmmCQG:WRnYT\gP_fOiVWc[
T9JDBoMUPOCi1oMUe:eVb`5fpCj6<I\OaMjU<lJISRP0=CF5n^1<dU2g^<NbZZ?I
STK>GTkE`L0Pm6bV3lgY3==bQRNnITneMUgn<F9q8BA8d_@@0Y_d[]bV[RIdV9:;
ea6Y14km\AV9WTU3jmbl2co>Ro<H]9iP8:R_mOAIQe90_=Ek]=0hp1m`ReSc7Ln7
0?feVoJ=1gA9]8ZT:=7CQk_ehljlOf[X__ZCfEGmFO@4FB5@9Hj`81KS<8lLJ?nE
@EB_7GgS9RKEP=In`JH3;6FLD^4qT;IXMD9RMGa<Oc1q@DTU::5fho[4N:]M38U4
ME0@SN90mKH2>MM<=AK`jJg9NL0ZXZYhL?i4WFE4TBfgFl1]Sg\>3UUPCjVp=I_9
3M0cAl3GclMKB^FQcOkA4A0gC4JQBYa16o=]V[UUM9ZZ1iDn2i8oFOjc\lYE9mNc
K44qZ:7EM`X21am67X`NIKSI0BWC47?N@LUA=heEM3jefWjEoZ6U4h[g6OXom>f`
O@39<2<MQGV0\NdLXX`aIKSI0BWC47?N@LUA=heEM3jeb7FJm0KlIV1Z4iVh?g5[
IG4h_YmcED^NqNSa]1R6Zmf5\dQROn3f8L_GJk[I6C03=4_Ec_mdjOd:h96@U^;n
bAFoIlY[6Z1fRYPCNTI;:b6<MSQRTn3f8L_GJk[I6C03=4_Ec_mdjeGH9ATCj?ka
U`6B@T^geBj8S3:h=Pf=`pT?;^m3G\<1ZkDb8n9f9AXik=:KcTZ7CB[T=YmbX]1h
<UoVYKJi8?h`>1:IBgJ:WTYhO7MEVJUXUn62Z^9f9AXik=:KcTZ7CB[T=YmbX]>k
:;i40_fKh`UPK^I5?7^gWB5hghM_e`pmY<5Cf?dj1dmIXIKY\ACUkX;1[28ZX9Nc
F5>j_2>c\1L9nI^P75b7<2Ao\I>j:0Wm8OO>ST=bL9[=aS?IWWVic^=Ac<iZX9Nc
F5>j_2>RAW:S59;0JR=8W59b@[`_?\X9`3RldSNp4^Glj7:1AAoKd5EBNd;2LXEL
::mhhgnNmYB?MeGd\IbS2[f]lLmT^>Zh>MX6Phiqfoee7oSH0;:>BPDdH5N88K8h
V]TEUR<R^0Vc9P6j_gL[IjOQMQJ1@\[VWRGQIB8=GWA2\X5;>Wmm]PDdH5N88K8h
V]TEUR<R^0Vc9P6jA`2kd8=ekJ1VB?JfoAUoN]A9@C]ZZ8kKqH4]J[a7q3@;K79`
Na]a7Yhhqo93A9H<XMhU\onp3CJ??R$
`endprotected
task reset_signal_task; begin 
  #(0.5);   rst_n=0;
	
	#(2.0);
	if((out_valid !== 0)||(out !== 3'b0)) begin
		$display("***********************************************");
		$display("*     		    ICLAB_FAIL      			*");
		$display("*output signal should be 0 after initial RESET at %t *",$time);
		$display("***********************************************");
		// repeat(2) @(negedge clk);
		$finish;
	end
	#(10);   rst_n=1;
	#(3);   release clk;
end endtask

