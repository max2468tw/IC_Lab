`ifdef RTL
	`timescale 1ns/1ps
	`include "CDC.v"
	`define CYCLE_TIME_clk1 10.1 
	`define CYCLE_TIME_clk2 2.5
	`define CYCLE_TIME_clk3 11.1
`endif
`ifdef GATE
	`timescale 1ns/1ps
	`include "CDC_SYN.v"
	`define CYCLE_TIME_clk1 10.1
	`define CYCLE_TIME_clk2 2.5
	`define CYCLE_TIME_clk3 11.1
`endif

module PATTERN(clk_1,clk_2,clk_3,rst_n,invalid,mode,recieved_data1,recieved_data2,message,outvalid,out
	
);

output reg clk_1,clk_2,clk_3;
output reg rst_n;
output reg invalid;
output reg [1:0]mode;
output reg [63:0] message;
output reg [71:0] recieved_data1;
output reg [6:0] recieved_data2;

input outvalid;
input[71:0] out;

`protected
>f<[4SQ:5DT^<12HdF]ci]RC]i>KOgl<oMSAoQ]9n^d_HUM5C1l4=8Z0RbMB7jWD
q`QA=Wi7Dh_?[2?kEnIUI:FX9CaUNBg>0aRhX3ZTqAhV[iT4B>E=XC^Ula@IU3J7
YUHae^895kmM_=Le4DR@]Y2Lj<[<SplmWT8Lp6[5<0c4\Dob?>2Wa`[n?6]^7O;Y
J:^5ngk`nF\b6`4:`a3LGV6p6?J<8EZY`E8eV;CGU;lG@_IiYK7dT4\REZV?_6H8
QPn1EiV`4mqOUb9?jY^]kPG8F:_<dU>Y;8d[Hd[l9Mb09nFKaPBWQ^?OQb5O7qO?
gbh<HLUlhj`O6F:TjV7mf]PDS[dgWMO@HbDi]2PLjkhQ>8o]Nd4VEQbIpJF=io[R
:9ZBNeKJ6?@5]Ri>WUBD_cm9A54a[?Ui?mTiAMX9\2X>?il?i><S6=LDZT<q==;k
YBEfMD\FmR8o62S6hWqX_YLEY?HE?1AQg?4Rk8OWcDcC5[2>c0Ue>VM^7p8H_aC=
9hCYG1:kn[5[biD9oqZZ@kQ<UHd;dQ6VFkS>mI6c`>BPeNo5V;gYDfRALicXqaZ<
;FlqJINdjXpjHe2YfQ<A\d7WV[7MSXNK@K^]1VPA>qhKdBC8^BkS0k`[H_FG8N5B
]NDX_@h4mq8f2OLZ7=>>AC10mebfO7cTq^P;lf=Wo`>\Hn5iNXXf=3FOCbRai[4J
[\hCMMigap3LgPFRh0E:0E2nkdJ4cQmJJa`803L[lec:qcdBN`1AO;iXfAC`g6F>
`6dC2Bf3nWDFLoWF3MUhpGXgkNh?oYhC7jl1gOOCPmT`9nO8TWQ9Q\>6QTZAoYbl
U\jo3WGUS__>fjb83VRXIj421A^M=9bq1oD:T`aHmNRkiiQGU_dmKkc1jCcNQAG_
E0>P68fVS8=MNj7phCma>dMcH4;WK_nMTnhGlaZQYKOOh]ccpVMTBS4pX`XD4OpR
aPSed_e2^jOca\YRcN2Y^D>FkNMKBP\bJj]RRJoS]AmCaCZIcfY;B:K_^ZA0D<4@
4SLN6qAEN0O1q8hj=RlplSDS<M;MVT[[n9:AYh:UMSIE5@V_0dASR1G@GW6cM=6;
R@f[RRCJ=IZ_jbGpmh9EX8W3^B0_O8mf@g^f@X=jQ`q=`bnO]0:N[STX=DU5SmCW
kh=JNh@4RcOLDaNAi8LmePODRhl:K9@BFPcHb\q4SPIc9Ef]<iC6fi]?bLhS0Cji
Jq>^hPc<OEINUiFSU_9n7jX=4?PLbOZoU:dmnl]1GESkke2gKT@I?HPc=_FK:qh<
U?TJVn7aC]Dm@Jl33OB;[FD9p?P56KdpP:nEg<9>Zok7]9aX4`kGMQB[_1Ee=Edk
Zc8e?GV1<B@\>G453f0lZh:jiKHE13;C=neKOeq]<?8UeE3T`q8@fG9]qa\<Z8I5
D0]KC26LEZ?V\2eAaWNqSEG[KgHhhSb?eNJjkWd7XVC\glh>[n:d\IpXZUN28L4_
ECLO\\3@j1>TN<DSdPAeeJCm4Kj>AbWRMCiphi=9kIoA:DRHhIk`6`j<aB@OgQR^
fRl:W53SE2O:g^6q6l>^:Q50j4ca@kNXaghB8ZacF9D]Dk2aI0Qp43D:=Ge[eb5;
:^MHoPn9i3\Vd_bQ7WRTd]QkL5Agdl3^5kpFLPC=9`]3Onc<1V>6m`lOFZHEfn:p
6jioZ\GpcXLXgOZ:8FV]I`?`52FXOCEbG75@_G1I0mkWJ;6J[MHH93cO^d5Wg<\8
gJ3ebXleB8[m@ha780X22aMJQ2?_j@DmD_5Db<^XSo[M;KBaXbUqloCLWN4`4hh_
7@]l3AmKKFH[Th0?lRiWRjb`maIk8[^?eM4OJG5n6NahE[2I=[TN<YWZMWRFI<Vo
Y>Si;K1lnhgB?eiUAbLTXRj7e1X13NdhT^q<2^[O0DlmjEm9:;Oo8kUZEbIoj3pD
J8d6>fgPi^l\U>UUnXlk1W7G=3pIL4FVDcHb8F06gVaE8g[eLeC_d`poH>P[gOp0
7\WSc5JoPKLE]20ciRV]kOG=_91YDZ]nc`8qM<cN6eRg6_YkjiRT[gMT4\4:Ym02
[21_:9Mm[iL;4aWYSJDjCQ0A3hI0<Qc1]AEpE4I:;=aHm?VJYVlg6F@@TP=lc=Re
WeG;p^lcGLBpeH6_SbDpOK`iPj`q:KO=eXVfgP=mRi\Lamj[fk@TOnNc?BTH@YPc
21mV>H6JVeP]F`XYJQ_fH<]A<^60G6D7]ULDT1JodD\TFe86q96M?]Vi?X>?cWg5
=Mk1O97h1BWljaS16;V`dgOXZ5O24i5B^F^`K4fXpCLgJGk0jCVp;Pnd]`RJL3Ym
k<PNf;_^RGCp1\[gnkedA;gDf2=4_@5jYlDCp:AaDOfJOjAa<eS1=@JV:iPh^3eC
DpS_h^;G43JGXi:bTmkMeWa<q8><0G>gkpnBEejn^q8Ra9H]_>1GNnl:XYQ7[GlD
H3Yo\ebZg>0Zg7[mUo:bW;?\bH3]a30TSLcSkJ^\9B?NU:2IG<h>3T1?@aOVhLcK
9E5oK\946TeUUiTW_<<PM=9UiCEjpIkL9j::]Y`p4OSDQ=YX?LlnFANS>5d]GHA1
NTe<?^q2Kk0hnYfZcF8oHBUE7eHh44QDSqiV]c[C@Agn3nmHI0BYYeXC5\dRG^q3
OegCB5IlTg2A;H87UL68h_p1g:oH^_?q]Uo\8kfq:`>QYV4`7fLKENX4`?e<F\da
kb3pD6iP^mbp4ZHGCoqMaU31VJgE1\^CBH0SEJ]dhR`<oQ2NL@@971P5=qM\<IY^
EF7@UbUc;OTI3oU^I^UkI^H_>DS_L=RV=QPX9hOfc8qWg_DQ;kni^IIc^bYfgcVD
e:jK?CnhTC;lG`qM3T>8gGpC0Ik>0FnENZ>NakI=E[pE@1]`;XBa>MB4:Jk=FM;V
M>\3Me7XiNGO9MbPdX\c[]HYI2l^k_`3U=mB^GhpWY`Cj]NLPHQM>NbR7IgP@DoR
L=Z^`P4kYPe9ejegi3k_GkbQg7EnT[Z@CS?p0kUGXNAI7^LW@oaqVaUDYQ>BHocE
nAXi716;I0\;[f<X`<]l<cOdlBINIm^0c66bFUKgh4iB2SZ0_5e;a97j6U>PHocE
nAXi716;I0\;[f<X`<]l<cOdlBINIm^0c66bFUKgh4iB2SZ0_5e;a97j6U>PHocE
nAXi716;I0\;[f<X`<]l<cOdlBINIm^0c66bFUKgh4iB2SZ0_5e;aDYe9Z5JHgTI
?5K;4I]Tp@W3:hl4O7\2DXNI<IZL^a>e3lWfi<PhI0nlG^b?d[Q8n9jT8?mh6W2V
g2Q=XDIda@jWOT\457\2DXNI<IZL^a>e3lWZ9gBU@ZnlT^b?d[Q8n9jT8?mh6W2V
g2Q=XDIda@jWOT\457\2DXNI<IZL^a>e3lWfi<PhI0nlG^b?d[Q8n9jT8?mh6W2V
g2Q=XDIda@l?0TZ82^:MI^7k\OFG5qeaOJNGo8lY6F3O0N?nRk8Uc>T9;4hJ^BVj
4N=I=cdL<1Wm_E4kZh27LRI2U[Jng=\@fKKhf<O^>eFP^VE]Be8SW2`Tbjh0^U\5
4U@4cl@In?W2IW`MA5M7AL@XUXa=J2e@>Hf:Chh^HClI0P?nRk8Uc>T9;4hJ^BVj
4N=I=cdL<1Wm_E4kZh27LRI2g\LnJoenN5f6G_J]8NGY2VkO:bqPZkQRSEQZj8nP
9a\6V40hB@i24lY3nIGH8h>0Q<[5]]1YYZe[C?IdlLTk=<c?k4WfTaR3^EOZj8nP
9a\6V40hB@i24lY3nIGH8h>0Q<[5]]1YYZe[C?IdlLTk=<c?k4WfTaR3^EOZj8nP
9a\6V40hB@i24lY3nIGH8h>0Q<[5]]1YYZe[C?IdlLTk=<c?k4WfbhOC<^aoiR=H
=[]gEZ6p3BbHXlq[i9BU6nqZ^CcS7?Ic[A<31qHD5m4=LTB1PQ;B1NWjpC3D[QO4
mpV`SUZCC;a?bb<1XPR8:hMhj]e?mo1SPXYhqEHE]2B8iHgBSOKKWVQqM080SoRA
E`aaf=c:GVEqB>cKCiB:RG>e3LlYQPApbTYT7J`@n=Ol?JWgBPIqhESEMWldJ9q;
HhW6kqojm:g9n9Y2iVDYfZ3CMj1Lo2dIA^5=XCPQfP261]4CqJR7CK2^iEQaM<dm
b\FAA?]lFbeIp^lTFkPTIj;S7kP[iXOU9RQAK52m6Aiiq?J>NJ@NP]mLN3ICao3=
E6K=MjD]pZoWCYjXpZPJ9@S`qQ`^3Daf>Y8P2idG_GQ3:I\I1fO]G4GBoD2pVXT8
B`\SdK6]CZ6D0[H3PA57mcQjNjH3?Ha4`hqY5Z\GJ=XR\2AF:ESH16^A9>THg1mC
N]`W8cFec3Al`H58_^B9k=IMX;llaRGpPVo;85WJSY>5aSMYFf@_a?Vegeb3E:bO
^QebIg052X;<ALLpO2QaS`4N^>YnH[8^hCk]0jjho3GbM<DA2ApffQJl9VG62PYk
IGQ]P;[loIZblV=LC]^hmHi>Uak<@l_QI2p0HG8LN3lpX@O;]GBl[A28^gY8=];U
afc0fA81YG_oOY6_E0@6F3qfXceCeRqUf`fY<_0WKgUTadOAhGPkQ^CL?Q8YO2lJ
3f<7HnMpgPjXO0Wqo`69ohMZf[bX^X3<FlRc4F6KNgPZq3d4QFGG<88l8Ub@fng6
ecE@Ml_N`53>;;EBYq0L3?O75>cThnHj>;ld6112a26Y<nHiZn_?[W[jJZ_?l=kn
::PK:<VSYJCnQC6ED4T]`MB0j?qal8OF>R^TX?_fAkT:YDKk8<@ZaAm?@lUJ:IJU
GOF@0hWLSB;hCM?jkfplgeGN^eJkhg;j>@0nI=_;?=m<[_LnoA=DHh:LTL4SVd2_
DS7J`Lo6FDqb=6Aac?4e;m36P[M]<<TBEPfq8bAg]VHpAU_BbKFGhDDA9OUnJ:[5
`A^ZJRDqIeaiVV1d92HAGHD7De`\^4p6XJI>fGW?E?n:l4BPQ[Kk^KRM\A3OVdl4
daE[`Q`28[c;RmpAFc;_dDdT@SX3cFjm8YY0TF[ca[R@o8^RkV[f<pU?G_6IA=:e
7_MD2I^dA:@d3dWJNJ9:Hd\G]:5Sq7F?Ej::Z\9\Z5XGU:[Y;i?Q104pK;JcU4dW
X>q;7^]k5`M_f0c[I8GaWOnFD6o=2_4m01`KlK;[dn2@i7AlTME;d_5Qoq]NjKKV
qka>Ab4nY2i0Lj:BUGQlOQ4FMOXDepNSJO9MnR_[6l=ZMa8cT59Ul_0X:=Xf7qYH
8h@4NLaghBN?a8o95Lik2_I`QpEGMWX[PVRi068@;8U8fEWUX3mYfiBY6pcQQ^kN
QqXnEG86hqHM>99cZJg6_VSdj19MWTX?l`:=RqFnUZ9^:0?GF8il=_Pa4l6_DSYn
Df484_<H_bIKqTJAj]SSmVceTEE>QjQ1o\0C;5RCT3UIm9JRG_Z7=@^?LZRlp0Xm
]FFDp^M^K6^=SSChklZ`YVBoQU60noLP0XH:5`IdEl=f\[A0:UZC1gVM2f[aI2j1
E_U^AG`9^Ml9dSBZ]p]3WAGDGpoA:j:Eg?XYk^fnW[WOBj:?Ad[ZGFNW<FKUUk0E
[GK1R`i:qDhVdB3YpnDaNgfg\:fo725mO_e129^VU4_98k9qi>eni<mf]VY]GaQA
c1B\`=beNjX_GQ8@DajPqhJm6m7OZ4?EZT0SnIQ^X\edFJ7mbMaMojAIFPQY>FQf
alYmIc_h6R1Cp_V>GUil8J198I?YS]:89=fL;=OeJb:0f9E?UIMiKVlYbkcOXIhn
BWJq7McHd9PF2`W:hXMRD5[:2_al6Q1=5S1S4\cE^@lBmCGho]URE::`k88q_Y]a
\a<pFZU[DEII5gEI2gGFUD61GZA=qNDUSZ\NqRd8:bbENnMHT@W89YYqMb81^oNK
da3d<=L[S40nL@Qn7?mqW_7Blj@XPl@VJP6mY_Chc>q\?eSX`biGjPNAAH5gO`M4
XVS5f^OjB_?SGG1;XqG^C[8EmO]1:ji>:RdKVEUOWNMf\1g0E09nN7QYp4MhJ7MK
lCR`8gCc5VA4ghagNm5pB[mmL43bERpQPgI?bq\kiVdB>;49[^55;MOOjYJ`XWCb
Hc<66G3U<\A<=f9GX\TXWKO^7IEUdJg9JU>7pjbZljB6[6fV>KEmgP\9en]Z@Mn:
YqVODAd97DaX>ch_CL4Y8Jm3l9^WLFg[ao5]\1d7poLFW<f_\nXDhR<i:T=b8Ok2
IphW03XNWqYBS^3>[jmn2D@b\S7<Qn2:VHlZ`CpnJCQAfEkq]JJn2FAH>?U6EiVL
b333Db9Z<OA9cC5TV@Pbjak;Ue]B=LE_o@:oZARCUMCDYlaC`^Nj9SSq\NGh;5M0
clMP[l3CS4IAS[_5B:aS^Zh;D<heSiLf=A9JcgjbK:GCjIM8k8XZa<39SPVCd31a
G6F5pIR]J=e`SFHT55JB9EYTEi8;>7ZV0cD3_VZP@<N0>``44[V<W?Q@6EF?J=ih
lG2N74@TdDWQqU6?4g@EpYc@2R1>6[k\n=QUNGn==75OBn6AWA>7YEIcgQTeMH5i
9qQCcY0AN5YEP\RDW?2G7W_ZF4=QiJeF2i\0@8B?K0;??bmbQ4J\mPc[`\3??16g
;q]1gem>:Pq@F]kh^>8C<0njKeN5?g3;aFdXO8Q4`V]3`pF:3;_eM9p9=c8n=[i;
?J`;L@2mXoIA=\CoU8[^hD_V[o9>JiPM\g`M_X`8[qeTcf^9Mg3bLBjZX5CPmK<m
[bQ>Ui5VQVGM_db92KROel5MSEZSqMef4Ol4_O8j`RW0cM[@EBnJ?[?_hKOF[eF^
kL^5Q4ZD?eaG\:gqomFaW:Am<?S<SVQKHjQ?XcBlm45IgcCA?iSYL=<HFCTjJ4Id
Lap;1L;Ynb\EKKcA?nb6Cg8ZGg6?GCfQO[i`@nXl[2bF^UFKI1X9LX;lKe`bAcWg
ko<CocjD6pHbRhm?eD\PX[ol^e[MXhGYkXNjkA=XWQ^66YT1P\h>nde`40<RpG;P
M@cRfO^\oW0_j>Ge`BDKej9QaW=PKUahR:\Qh`eG=ZXRKB?q<ZJob`SAWc;X9SZV
CG\46k]deXMTaelAH]0Nd5@0>^3Q_=VSkBq1Q6E2GDL^eRd4Um?QiCTG\nNY<n`:
^k3Q`FR3^\G4U@=RIQD:6q8Z;CYb[TV97MV^iPYBfdRdGc1N<59S@@m:0=X0Jcbb
]F<_goj:po_aWaO74]8<E0A3d40LS2biE`o5[2_fHR01Kp<XH9N4JpZcoWTk7QiB
Rk4bK2FFWH;]T@7VVMKi7^`^S>GV2iOPcKp>LW;FifnNkWf>^KMbM5g>nPM4QQT\
TfjeGdI=^2JO>LTpT61W@H]>eJj1S77B:T16:H<YZ_PlEA@E\YGlSIcnG<d9pEbP
IC2RRXQjV4UE8JRj3_PkE]JK[4@\^ZcJ:_OXhWe3TqaG2IRZOF<_g:MU7HeQXn@W
jkf_a5RQ=3:?@SH2h?RNEG:51:0@a^Fd1X=^p[[U76;faN]>`?Z>UOImm?E7CZeS
LNf7[d[@T;Y0:ioVLqo3@8U>_IT\h\iDlEFOUUG3A10m^nPNekmKAT]jKoSCjcp4
\S]C9K=EPNh6X>>1]\6D=bAJP5YRc_R1@f^?F\Xg2i]q]`9PJ_8H9n`XkQgfkdG0
9BAIEM3dYE;96C[b@Uime1I1p;VQME?QfFPYl`=bNm\9Y@FmocbRcBhX9KA5O3c@
_p]2CYkT1AaUPX[J2=PQ0Ipg@cf6D4_@BH6mDd=:1ZYeZdjJSgQ=f3P3<;;V]A]K
4<noIcOVC[GO:mh_REeM27pKcHWTmYqOWZmKYWBp4lZA40PqJV1ZEFhDp>LSA9ZC
_pGRHjC487MndPRAoZ`gJC=W24<2T\oj=3`>BRedKk]0]1qZR4Ql]A:UXBK9QjSV
KAQ1ZP4C1bOpaag<M=eT2bQH_7n0LRDHFLUQf^WX>7D2;lo1DPK;Sm\Np`DF4a=M
M?dI>GIaR_ZWTCdLUE4QBIg2]:h3P2ShEA5h1p9oU@4_:f23]7V>SFLFTo`MR=i[
`7cl5i>hVKNieK6Q@oqH7d4U4Y?U1_AO`QV6WC1A^?@c?BjPRb;n?e;I2XQ9Xeiq
E?o@TR@8am>a9]7[ABSV\J[70FIITR@6@9JG62okcJfQg5CI2YEAkVPgF=9KS=p_
di[Kfl`BlP[lnYcPE;<O`A0SJ>R>naFP;UaO2]aPbNRpaf5:;7ViX[GMMQG14[5=
nP6HMg:iaMgCTf<VZX?51eV^q0Zh?eZdXj1BMkb_c?LKU>>G[\MeWC:Rn?RhSA_D
0F]l@qbLfPVB`LQ5Dl`WKMR]aGpX6PmD3gQHf5;bWo;K6D`ZlFO<?LTe]GTV>:9m
HIH6LEcIaA4jI?W0[NUPTNI9k6qjL5neTJqHUIMcIjW5j=B4:gI^GRgCNGUpTPW[
SDmPp]`3j6`Xq_8mU;blfqbVM9GGOCGQBUDbEClWYVnBl94aRl^?6AiE?<cNM2^b
4;TO]CqY8QVb@V3cZX8ia[d5L_CDPaN<:@jO5EhjB0g0ERX;5c\IG@@KhG@ZVS0W
9`qN_N1fb^E6C^FOF9Q2P0J6PLB`:Hah2`51=^FbCJU<1TK8=jmaD]qQ^Hl:;7q5
02hLQmQq]H_1n7Gp[e`>jjgeHnPg7E<e>b0oL8[RmhA=DnViRGBbQV4>[QhV6^SJ
5QWg3PDYXL8AAT3[fBB7:1q9TV87cm:q37X;Gh^?qIa`fedh9@Gh^c=C9D[;A@H`
I06`Yc^DFBQM2Wn6fl[I93d\E^i1]0dV[H5Mg]amYe`1Gij^DqM[8Z<FS\5]Pn3I
jRbmj0SkAXTMhJ8G<k_08Bjl\5RjmdqIkH17WhhpnmH[hTI8D4hXiVqQD9g91JKa
?hCZ50H\ViEF_CW2JR[aCXFlWpa91S1Wm`qU5iQIHM?SJa=<l>Vcncgb2l04?:NR
oR0HVBU:W;L^JNO:JHkH8pcZBFS>O_WbC6=B86MYPe8=O2kdN5TVI=DeJTOk;O\T
m`R;nk?=qd\3`g?HfjEhnToY2T4A<CjRXPH1foIPCZnHgZi?FiAGT^>?7@>pjHe2
CNn5CCJge[@<]:^Y2m;W0Ob?\AlUa1Q5K8<ab_TJLlg_?VqFjmn7Xc;f92MIAgfA
JR4jI620AB3CVG@o^V\KO?Ubg6S1c1`C<qm;_k9;2>]fIj;OX4K]M]o=jLd[DDj5
lXG@MJ=MTKe]in@AkU0>q?Z61:j\nh;Kc0=eE[O1R?hMl9JV;^nmCi]bZ;LIDem4
FGhbd3nqlAaebK5YdK\_jG7pXT?U6oK;_f5:JdZBVYUk9DeT@`6BM_@Jm\IYoABH
idIWBR6F45p`UDQ\L9FGW]8O[LPY7\ZcD^;C9HLZc_cm\7ODLBh?Q]MGP^9\5q;Y
P>3JipDV_YlcanPNKcOMGgnVeddLK=kSYLO[dJ_m93V6Y8TkIiphFoDP]B4LLJl9
m=Y=\0n0ea6[QJQMe9KSA26TW@6IQHMql]bh<3en54Zb`Q;jiCd?oPWBd4NWSMHc
M22Zk\<Cn85;qBEFbj>8Gc?33QPA@LJDVVJUKA0Km<]>1:jDaIWUfS=X5qX]<YIJ
U[^=<[\NMJ;7Of@A<95dZZ_0JN8=HbH>3jTleDqOCEeA[Ge`LLcmN50gDJ:OD82M
ldCg6VEheIW6^F@[PA]qn3eQe<o7W>giNmm]Uce9Q7;M=8_RXFjWVTX7WNV1DgM8
5S2QFjlmNl2qdBXP0R]h5W2P:9Da;X:l:cnfO72BHDJ_@SF[acg?]PP<pZXk4N:e
PiZJoGj7\?LGP>ZkoOHM0IToh8?G>Y0n0c;M[pXkRj7YKg74ge:?H<<?VKqUnH4e
8i4GkRDn2`dSdd=m2;^6`COZR5dYI3XPc\5[aXblEFW@K^U?WPJWDO3jM5Vq5fQQ
XASq@G>9T7\iqd8939NKqYbJaDh>\O@@7QbD=n;XlDmkK0UAN5Z>YE5c]1QMZ:bZ
Lf8=cYQ3WcolLO<`JSh^p62kKU9i[q7JN\T6O5pJ[5SBAgDEn137A^Nni;XmSjH;
eMN]]HZiU8:@?\RI0>nqE><\S92?_aD;0?Rhe>GifOlVnXlV[=EU3URSBo_IMfDi
qlD5j3=h>ePK`QWl9beJN:R8i:9J0;f:2egfEbo9dCFmPpMm=dMGFJig5Pg9L1KN
F]fV57A_PR4lj5:WX1a\mCn6=@qg;TPQSF[24O;8VA?@;=1;J]];nC<k1B0=87Ne
FD38Ga5pk2BEZSV1=:`6?[UV`^D7UX6GBhYFF[KB;KOj\<mGAbS^nXQ\F;bmcEl^
nPP78o4]0?>pTBf@OUaJ;cbkYoQdfK7mN9?X7GU]]]aUR?20>aRCShk\qbPQBSag
`TbFPZJLo@BJ5M:S2;Z;VPDdA7CZVH`Fb[h\nq^VWVVVNe0gU1=hbB`0mHjBc\bf
Dk9M@8CC^kmIm\G<F^qCKoI6l]ZLJi]lPE[B^cepK8R:18K?kdaMg\L2^RF<_@_=
b`Hj?;:U<f4Lo:jgTkKebG?BUBh9bKd_GdfVZnD\qQVDT4;1pB``m\h55pSa\eNm
<p3^CA0Q?\gBIHindDkNXhHCUP\1o^Il<HB`X:K\lpaCKK`_kIF;?Yo>j0`epWaV
]DjHm_@aLJ<DI:UDEq:knJogK=Z1q3k=I`[MM6e1CDSc?U2V[T\qF1RGh3nhq;Pd
;\ZYq2gdKeYX7qJaMY6YTJ?a0e6gAL@=F;4L40>K9`af2OF9OMmNUSC]\\QZ\ReB
:1ETPHYBHkc3Neq;oVHGJ3qSM2GEAIqU`mcfojqKc0WLe`5Qiq1W6Yinpcb63g=4
jfl?QkGk>njndXi0ZW]g<keL?pHJoOMF]4gHoW<f5b<B7b0ARqXFGO:FY]9c0?J<
T]`PSL=Hfhjfcf<miaKBToZh^_2I?0jZQYImLRHCg8mD4?Q2Lnq3KDHHoW8RZMcc
h=_FgZE\7E8F=lp3nmG=iXC07J[AV=ohOLmXT_7[?cW1Giqj3ZH6aiGjENl1f0lB
OTHf4RAOHoV:MqMCijHcKoG=F<D3_pkh86G5CRiY_a`lN9d]:jeaWkBN_m0BLAm@
PA`9DHY^M0:m@LRPFgf765Gk_KPjFD3Lc:>_CmiY_a`lN9d]:jeaWkBN_m0BLAm@
PA`9DHY^M0:m@LRPFgf765Gk_KPjFD3Lc:>_CmiY_a`lN9d]:jeaWkBN_m0BLAm@
PA`9DHY^M0:m@LRPFgf765Gk_KPjFD3lhgdD2;fIAdDJOnUcDiqm6@7G5AIWUf[2
bR51LnVgGR56bGKUTWm3e0I2;N]QXD`X;GHY8A?f\@XVNgP9WCcmf6D;hAKWUf[2
bR51LnVgGR56bP:dD]<ie0B2;N]QXD`X;GHY8A?f\@XVNgP9WCcmf6D;hAKWUf[2
bR51LnVgGR56bGKUTWm3e0I2;N]QXD`X;GHY8A?f\@XVNgP9WCcm0R>;Rn8c5TJG
j67Mc>EpB2AlRL:HZdJ4=3OU9gg=DmLN@kB;;bNQNP`=S:STmJoOXE3K<Xl8Y=5>
?EdRD=eUBTBeIG[a6dJ`=hH@NgYQ>KS:@hI4<b38n2o:DLVhm5aYkifN<\]_H=ba
<idFD=eUB\2Z?G:0ZdJ4=3OU9gg=DmLN@kB;;bNQNP`=S:STmJoOXE3K<Xl8Y=5>
?EdRD=eUBQS_?>>6lg4SKRQPiGfTpXP=]i8[SinADlVJA1SQ;ED6?hDe`GfV6Yd8
G\VY2_lDm<dLj=K:Qj;;`fTd7A<=mVf^n:V[_inADlVJA1SQ;ED6?hDe`GfV6Yd8
G\VY2_lDm<dLj=K:Qj;;`fTd7A<=mVf^n:V[_inADlVJA1SQ;ED6?hDe`GfV6Yd8
G\VY2_lDm<dLj=K:Qj;;`fTd7A<=mV3J]HSSG=N54830NDM=QpQ<^4Q?qn21\9EI
]jjGMT=4TQ8ojfXHlmZFH`B;<CfGgMCb[IGimG^`ifki>[]3^W?XgI7iqG:GUC4\
@;Tj9iJ\>HeNa>SceG7:OI\Rq\5^RkBRRIU3@0jN7^[qXmTL7_cUp2?1^WW2MJR[
HKJNQL>c>CeCpVM=TnZd1qFfK_Dn<M7^h@2Y0LUOc_OKQI]\Lac:_kBEk`\>=Jfj
D502FhV1oY83]aH\Xp9=m@eWe7=ap>8Y6[fQWN>>UC]QC<YIm<cYXffSI^R06XjJ
h0`4E^_O\@fXe^hjl>2<YEJ=RWcf`87mp0VW6a<p@@f`ePDdcZfK3LK=;nEg>0k2
5GqS>87L1o4k`JSSoLmqLL8;GI<Y6V]5JY\@n4IUW@2pPI9mJ<6^pXE^7CB?_E;7
9DiSB[cAqJ^Qf<:l;qgVF8k6]ZJ0I_c5pAW@dgRf@:BjZ;A`qd3TK8QoPF=4c0^R
2AAMcKch_8@?fQV17=lQhbm]\@QgeTOVTA>KYIl5?b`QXcV7e@@HHUeo>F=4c0^R
2AAMcKch_8@?fQV17=lQhbm]\@QgeTOVTA>KYIl5?b`QXcV7e@@HHUeo>F=4c0^R
2AAMcKch_8@?fQV17=lQhbm]\@QgeTOVTA>KYIl5?b`QXcV7e@=b3JALnEPGZcZC
00R=fpm@jB;>fRfB\OIlNjY=?koMS8SoPPfHH^4ojO]a:GL]PhTm?[hV_i88NDNN
0TXS2]mMjgDhfnfB\OIlNjY=?koMS8SoYf1`L;1ojh]a:GL]PhTm?[hV_i88NDNN
0TXS2]mMjgDhfnfB\OIlNjY=?koMS8SoPPfHH^4ojO]a:GL]PhTm?[hV_i88NDNN
0TXS2]mHU@D^jI66dhA:>heXk6pFgo[_M>FVl`n7fQNc?>A0Z9d9YO@TJm<Y:@8Y
BDPl7QZ;RX:^SLem\ZY3L3<2\:fFmD^QW>7Vl0NiTbkG2>1gZURAg1GTENID7@8V
hDaJ6gF38blW9Lom\ZY3L3<2\:fFmD^QW>7Vl`n7fQNc?>A0Z9d9YO@TJm<Y:@8Y
BDPl7QZ;RX:^SLem\ZY3L3<2\:fFjGEQ<dV`T0GfNUof3m5q53mWJTXaP7TWC2gb
mcTWS^]JQQUhXTJecjBg1=gia8cj=>6ddhh2]^NOg;gC@4X;hOof>dXlP7TWC2gb
mcTWS^]JQQUhXTJecjBg1=gia8cj=>6ddhh2]^NOg;gC@4X;hOof>dXlP7TWC2gb
mcTWS^]JQQUhXTJecjBg1=gia8cj=>6ddhh2]^NOg;gC@4X;hN;hHL2DXWT=3U_=
_g?fpc>ReZ\^QDF?]eQIb9fAGKCkRN9]okZ`FWAI@a0\gHUfU=9kUW`C8g`Q4;_n
kqgM7QK5G1O=VLY;gY@Jm5RcN?7Uo9E0gWp6P]0fciVV5dRSM1JA:plC\k2[NeQ`
qmHO0]J:pUmh[[10f`bJ:cJG^aC@]_GaXqHl1T=;^jpOJlA_Kg6:o8RQbPq_CJ`Y
]e^CMIQcFo:Hmf6U2U81@L[3j86072V5VV9c76?XPZl9=RhZH4B7=neFB0?p;n<S
KON3ZdLnNVV<ojmLBF41Ce]^[f@Xe;Y89e7_9F_mFKghE6@i^76k>no]9;hMjN22
FiNGZdLnNVV<ojmLBF41Ce]^[f@Xe;Y89e7_9F_mFKghE6@i^76k>no]9;hMjN22
FiNGZdLnNVV<ojmLBF41Ce]^[f@Xe;Y89e7_9F_mFKghE6@i^76k>no]9;hMjiXj
l;oWmK`I<bLn>\RZpdBaBL`YbLMgSTZ9NePXYkB^1ldo6fQDD6T?LSNmcX>JcNm1
ET@^NK7NV0Tn4l41<dh=ZSmY@LMgSTZ9NePXYkB^1ld06<j]NnT?FSNmcX>JcNm1
ET@^NK7NV0Tn4l41<dh=ZSmY@LMgSTZ9NePXYkB^1ldo6fQDD6T?LSNmcX>JcNm1
ET@^NK7NV0Tn4l41<dFkKSng4d1:MPGIclnS`p?>l16YMilk_7G=k<1f2Nlk@eMm
SS:jADV=8L[6SX3H31^__UR0Ih^bnac6J2Pb=mHTlWTZjoX\01X[cKTnHonk@dMm
SS:jADV=8L[6SX3H31^__UR0Ih^bnac6J2nN^[?d`?^_D:P80iDdmmnZS[lk@eMm
SS:jADV=8L[6SX3H31^_\UL0on]?J3k<UWob>dFmpCXoiHHmDA<;T;P>RFK5b\B8
GY5Y]4d7OS1?2;V>kgN5QHKhD_:FPIcNkA1@HBSnhCR2nhcnjK`=1X?Tj0giWLXM
e>hEcTQ7ITB?X;]lWgV5Q`f213@_gI>_ei\@2BoBhVRF1d=IZK`=1X?Tj0giWLXM
e>hicEd7NS1?2;V>kgN5QHKhD_:FPIcNkA1@HBSnhCR2nhcnjK`=1X?g0:gBkAB2
Y^nb5GPGh1PqUbAgST^Bmg4Ll>o_h<`7@dFLFoH;aMHH7ND7[XbcnA]GkEEYS6PS
dX8:;IOKhd>]oFVD0Y^Tmg4Ll>o_h<`7@dFLFoH;aMHH7ND7[XbcnA]GkEEYS6PS
dX8:;IOKhd>]oFVD0Y^Tmg4Ll>o_h<`7@dFLFoH;aMHH7ND7[XbcnA]GkEEYS6PS
dX8:;IOKhd>]o2LW;RTm;DRW[Kj_NdE9pm^47>0fIiR^<gD1WYoUL3LN]14^6_\T
6IKpNdj@B@P7U[jegMP\?jL7JfkL9LoEgTFkpbKdbG=nP:]gF5n9O6:q[Y]1b2Fm
pg_J=eK=UnHF[hnfdn\hbg6dOpnl<1>EeZk4=YBk2TI:UJpoFhO=Wj8FQpZ\06nn
;q_VZI`^bIfBR1LiGSAkX2L23HM:CB<ii5=<[TplWI5O]hqfoR]lTOeTBp=_R;l1
keSO?l7HCeVdgn<<mQ;_`q^9HIA<V<HcoEP23KpU3QCGFXMD8CNV\V0A\OSm`3p=
1AIAi:XqnY<kCP>;go<@If3EEIgqHUl6\1_bqD?QMNm>eV@36Z?3p9biPoi3g@=C
=ZfIY7hHa<:e8o?3AFabSO;f78?>Tna8eh[da=_g6MIapSEd760f[Q0<WLS[Q\Ah
WS2gk`QcjjfM4Ed^DlH<>0MIjmX0^>=?heR\Ej=6M@LDF_eQW8:fdQ0<WLS[Q\Ah
WS2gk`QcjjfM4Ed^DlH<>0MIjmX0^>=?heR\Ej=6M@LDF_eQW8:fdQ0<WLS[Q\Ah
WS2gk`QcjjfM4Ed^DlH<>0MIjmX0^>=?heR\Ej=6M@LDF_Lo2iYQS=o;o9BDA?XZ
Wpc3UF[Bbj3N3Oac^CUTcKoCZf8__0PAnYB]XVci<I8N[n\=]mZ1K`LogXXm?EQZ
FZcGRm=>b=3N3Oac^CUTcKoCZf8_<1`\W^c]XLci<I8N[n\=]mZ1K`LogXXm?EQZ
FZcGRm=>b=3N3Oac^CUTcKoCZf8__0PAnYB]XVci<I8N[n\=]mZ1K`LogXXm?EQZ
FZc0d^=RAjNQ7\mj3BQTjCpi5C^lIQ0Xa66XhaBJURCkE8?X@J]:5SgIN>4^`aKM
0>F8=3>0UF8g5?0Jo=jehIYiW:JCGQhXa1c[A@HLaRMUEMD]TA?:38BA3>BkUa@g
i?9;7d_iUF5g5?0Jo=jehIYiW:JCGQhXa66XhaBJURCkE8?X@J]:5SgIN>4^`aKM
0>F8=3>0UF8g5?0Jo=jehIYia2nCB^Wbj1c]>LdT3Ndq[@cXcO9kUZYI@B7Da\NT
ARMU4d:`cf`4P=]40CTS?nRK`BZ\laYT3Vo`f54k`7?T=me\2n9kUZYI@B7Da\NT
ARMU4d:`cf`4P=]40CTS?nRK`BZ\laYT3Vo`f54k`7?T=me\2n9kUZYI@B7Da\NT
ARMU4d:`cf`4P=]40CTS?nRK`BZ\laYT3Vo`f54k`7?T=LBA2SN3Nf7g^1gh@bZh
qGmjOXJh[W18D<IK]ZTfXW1d=1WZfS<FNq0ak7f13IG>oRoZ[K:1pZcN\0[0^ZGp
NmRS;^8f`K@2D8W;MnUeOb0SE`kWAVQTcAAZj=PFbXmXbY_FoXB@HVmaBkQaq6nZ
h7LhmalANiJY>aYF@f8<hE8olE@>WgA^RYVYIMSUHpS5Z4LhH4`SE9fM[YbZ2XFl
kP8kpOOBWF712pW_;3QYS<2QfeJQ2pofdKn^Dn7dUhj5G9X?7CQ?f7K:^8^Q5ohR
kjW;e36`7di>nbQdWCJG31=DKmf:\68VL=5KDU7dUhj5G9X?7CQ?f7K:^8^Q5ohR
kjW;e36`7di>nbQdWCJG31=DKmf:\68VL=5KDU7dUhj5G9X?7CQ?f7K:^8^Q5ohR
kjW;e36`7di>nbQdWCJG31=DKmf:\68P]<2@li[cE[ZHI\?DcRpPXaGDdDlM>2^h
kR[idDo1>b0E^EP`o`e2lFa5`=f:Y]?RVHO3MMQMkk;V>3f:?96PWM5H>DQM>2^h
kR[idDo1>b0E^S9TVj6;Pdn5`=Z:Y]?RVHO3MMQMkk;V>3f:?96PWM5H>DQM>2^h
kR[idDo1>b0E^EP`o`e2lFa5`=f:Y]?RVHO3MMQMkk;V>3f:?96PWM5HHfeMS?>T
DZ5k6_[@G<:q]M7Lj\6;JDZ=aKlAQdPi14K8^:`M_`JlJ1K9I:I=QHKdVHSo3Me@
\EoZ?l`=E06;:IVj^3YlJISA95jK1b\kC4K8^:`M_`JlJ1K9I:I=QHKdVHSo3Me@
\EoZ?l`=JegU]`4M7ZMP3DSCHHc1Jc`K14K8^:`M_`JlJ1K9I:I=QHKdVH4;DMQD
3d<]QObi90MaE0pdb[g1e_AQafKQ<[OR;Q8GNK]=0i7cmfeL`gYIg_k3K>5PVC6X
>31ZSUdHOSYbHL_dk7I2V@4fUTZ`W<YE4SkGFIUnMkB\c53Lo:?IgPXVKPPPSlLE
P4nhS8bb`iVbHB_4[7I[SaVjUTZ`W<YE4SkGFIUnMkBnJfeL`gYIg_k3K>5PVC6X
>31ZSUdHOSYbHL_dk7I2V@4fUTZ`W<Y8KS>:nKdhc=dhRcmjiVqVF^]@N3^5P_OV
EDE@UHM3H4K0LhDXaY0a1U?ZfPG@1_^VBJ0VPREIg1?h:GqF`F:2NgHb[<55hUTn
;U6WfXmVjYnH[9>[Xkl2d?3IKlW5^9ESW\RLkEVPG`5[CM?Ki`g>Wg3b[<55hUTn
;U6WfXmVjYnH[9>[Xkl2d?3IKlW5^9ESW\RLkEVPG`5[CM?Ki`g>Wg3b[<55hUTn
;U6WfXmVjYnH[9>[Xkl2d?3IKlW5^9ESW\RLkEVPG`5[CM?K9J1a84XOj6^PUgH<
m>_pDF5E?FMV2B>cNhJk1mf\VgFn26_@oJ5Qp3AC6\\_Va5nXN3c;oKq>cn<L2fB
q63TMd>Blge0e:KjiFl0<5NeFq6[24QdXeQ3kYiG\_9=5UqDOUn]Fe4aoN>F0R;P
i_gTGd_T^SJ3S_bhdWCH\2K4Y1OqaH:i20PfE:p0:nDS:2pWakcHDep@7f0gR:=1
HqFFIf::_6C]_YIYk70<EnYeM]F39Wq91ImG<E_[CoXAj>adaNdK86FA=[KP^q?<
e;<1TjNZ`i1HSXV?W>g;j9[<4GFl4cS41Ne=6faR>QDLD7FljiI\dPYjjDMU]3PO
WP\NTSNZ`i1HSXV?W>g;j9[<4GFl4cSV1^KKRYf11>2LD7FljiI\dPYjjDMU]3PO
WP\NTSNZ`i1HSXV?W>g;j9[<4GFl4cSV1^X9TSjl_lH\aZLYggp0G_7BT3kgJF1d
I=j`K4OHWDDV>JM_Ndlng4^`K;mBDd<aJ7TcoJbh9Io0N```a@2^BI9a83XgJF1d
I=j`K4OHWDDVMOS:eZN\jSLN^@IVL@WS6EoGVJRh9Io0N```a@2^BI9a83XgJF1d
I=j`K4OHWDDVMOS:eZN\jSLQD[]L9:D2U3Fk:Ffq@mLeDeHD1K;\o35adNm\hXUA
gcK]GfJ0F@ke>S7A7G0hmnQ@V09=940`iXJRjcZI?OMf20HH1K;\o35adNm\hXZf
=dI8\TU9LOmNhBleUJBO];Z_a>WLK10fiXJRjcZI?OMf20HH1K;\o35adNm\hXZf
=dI8\TU9LOmN;iDPiX2=MJcQPL]TpXGf38OEkOl41IT:i=>PS:?1G_=^Dcf]1WZ\
EULB^3ii[eG08c:HW9J>8KK]_ZiTo=i8ddaEhOl41IT:i=>d`hgo\46c@3<l]c38
\___4aYGj=TH9J>QQAbfOKK]_ZiTo=i8ddaEhOl41IT:i=>d`hgo\46c@3<l]c38
\_J6kN=U<5VR<g;Zbq0?Y5KVj6P1FQA?9Wena7VW\2NF^fEe5<R;C8;6Ad\aggW7
]:aeUBYfQHi36g8`G5UnhJ4IjaP1FQA?9WC0m[LQiE4C<@KGICKRHWYkGWJV5CHg
O]34NL_2:Yi36g8`G5UnhJ4IjaP1FQA?9WC0m[LQiE4C<@KGICKRHW:Y1[VLI_DZ
<Hck@nq_1TI?]_A]U1W<X_VH;WJUORaC<OSe\7Ain2Wb]^AG[Hi:TCpn>bD]?dWD
B=;X<iZOIOKhd>]oFVD0Y^Tmg4Ll>o_h<`7@dFLFoH;aMHHDEXCTfc\TLan08`\g
n_OlACCNYARYCCkJW7P;VUaG5EWeTN[`E9[:>g7T1alGDFCDEXCTfc\TLanP8`\[
_nQX<iZ@jC93\CkJW7P;VUaG5EWRhE]:0a3jKdZECjAp>;nVXZ;DVaLG`;eGJbBB
oNK[`2AT]KW`ec4QjS4m3P@L]7]QeNIhVgF2O<iG9g5Z>Y2>k?NTO@Jg[oUBJbBB
oNK[`2AT4oY^8;R7^cWoTKER<95ibURfY`7OXYm]o2DJkY2^k?NTO@Jg[oo2=3Y^
b_gO\S@LJZePK@][J5oeJ07N_T]IMe[kpFfK_\MneU<EQ3J:LY15]RWSJce>?=3U
7Bok`QDFNOYm73b?b=iNDAg]I<b<KJC@:FA4FZ6U>hdf:\i4[?CFJfjSNce>?=3U
7Bok`Q;1[;RklX4iJd<IAJaK[lLHSIC@fFA4FZJE]l^>223T4Y15]RPI5UW5N4X4
VcAQ3PV6`O9geBUcFl0Ynp=5T@TT1QObRFO7IA2O4:8k42bcL\1WY8D:a`^MX]a\
>[`XkNCT1PPG6Q7dn2k[dCNAABVT1@ObRFO\>EhCg0d4ZAH`NTWAAH^naV^MX]a\
>[`ggE2bKZX4^G8FMmXj6G=k5b;RW3WV5b9eXh2O4:8k42WYNMcGEFU<:HE^@7Hc
30nEL7L:@>phnDeSh^L17CPJWSYVKWNO9lboH=P^\A5E=;Jhkd>oEeWDXk_5[?ii
Xj2PND4l<G]CRT:S4^D17CPJW9?klc1lPh8cEVb37N<gUFX7XOG7Qe`DXk_5Udk^
Xjm0WJ5]Sdgh?HKF^LIa;ARjZHTVKWNO9lboHO237N<gUFXYQn]\b]67YjGQT?4p
9J9M5hImRT_>PQLj_bf@MUCBG9>;iC[2m5WhO_;dDC7XUIkBX7ijhEPA]:a:YK_G
aWZ4oEIJRT_>PQ3jOQ2[<hn<_g4H9DSP`kXN\5JGKR70]I;WEhjb@EhiDF[H5f;T
9Yc9X@i>V^MkEPbi_bf@MUCBG9>;6DS>`kXNAnbk\TTKU3Kin;YMpWIB=Sj_C2_S
E<@EB]kA<DPFI0cUO_mSD]JdNfapNZdWD28CVR4i8YjU8dXSYTo6\RAYINa]djKh
YXBMPIF5AT4D3O@fD92gkDkZLUemWib[3G8<lR408YjUA>e9gU4fP5^S8\0alKY?
SnDh7gG\9b8H1>QED92gkDkZ3D9_NVO?>Lf<8V_:hA5TcdX>YTo6\RAYIa0alKY?
`?6nP;6o8>RL4=TEqTTVFfYjA5Q7naZWlQcP?SDY:A>fRmA3jkm0kK9ZM^7eVmeo
ZAM<i;]NJVUj54CFOi@Pg45jA5Q7naZWlQnA80QVVU3FZV0^?89>;[[ViYff0U1a
CjKI8<oNaVUj54Q:JT7?gQb>_Pd9HQbD1lRbZSDY:A>fRmLiD89>;<\=I?FVR58i
gc`6fp3Q5;h<0lXLgYg;0FT6IhC]M]k`5_2Z65T=[RS>ViE44<@^44i`;h6QaBWo
4Xk0Nc]@Jeka0bXLgYg;0FT6IhCV2_C<]ElSl?U=[N8^Yii6_GWjOGeFRhHi2eEB
4kk6hI3VT>0L_l4;TDS?KiW][Sa;MGk`5_2ZW5G]62mZ8Sd3DRQleSDD2PpIm=R7
aQ:[1A\]?_mMj9JU=onAIP]mdTd\h4IW?E@lkQ:0U^7IM;8RFeOP76D]<KlAkmI=
TQV[1A\]?_mMj9JU=9nUO`NYdT01mX@@kEHlkQ:46AnYU7j_foEiHSRREdjIH^F@
lPhVMgPIDbRC;6Cl_T1^IPTmdD:E?H?]LgBZ;f=NXo\W<c@p]QJP<I=JJA1a0Yo>
Ei^Xl[>JGT:Se\Vh`H`JhBKY[<Je>7RSQUYR43L>RJU_dTV[LomRNT=cJA1a0Y[]
Ei^Xl[3JLU=8c3?^FT1mTBK[[<Je>T?[NcmgUcT57D\:?EPG]anm1JaXKgCm1K=4
GJ7hDdC^hT:ne30\CH`W7nFPFnJ1\@m2@o6npcb5GOF\2O8K<@\ojh1IXh1=i85Y
SL1APf>CHNiko[;eilZSj>8U=n1YA<S_de:c?_Q[k[9\Hg8K3@\ojh1IXh:Tk@_8
LG2_bidNPNiko[;eilZSjaf]`^YG`5MNe>acFUPCaSVRF:=LjOl_mAIRi:m=485Y
SG2QPf>\O_aP?DM1@WC9kX]iVq4;2;cJ@cT6<GYfkE48H:Jf>Y;fED5SQF39LS>4
ER^glX@M0i@D`MdCS7O]5;U?Q7QYbeXd@aT6<GYfkE48H:SJQ@PcECMYF]RaP9>4
ER^glX@M0i@D\A:I71hB==U?Q7Qh\]^SBm7=6Sal8N0<K\gN>`;f[AMhQf39^F1G
BI[W95`C4PJ0@^p]ZC9C:a?=@khVWMV:o8lehGFBR_[k?`2O[bdONVko[_>3`E;3
`pH387WkQm:VEYLBMdjX13PS<U9o_4;c@4XnF3iNMNVk\kME\2]JKGRh[ThMZ]YX
If:i]AVYQA:VEYLBMdjX5ZgV7e;oS=E4>QgWASFPMlVk\kME\2]JKG];=n2MZAYX
If:i=aHORD]JJ;<c6cl`<SPS<Un=5_;c@4XnF3;b>XT7eWKWSTD^Vjq_IPgbk\O0
kjlA;5X^L<Tm64Z2BghF5PCYVbV<Zb`j<ZX8?QFJe_IoYiQ5j5AKG`=mUF;F2]>2
YjmA;5XG^81`S5Q2BbZ=]NZ_LFET_O;l<ZF8?QFJe_II0>I5j5AKG`=mUF;T2:[`
3Y9KKo[__<3m6ENh8g3F5PCYVbVj150:3:FK^kW>ohMpak<mQQn;7kg287_5F^DL
UBfVL@_nPWWgFOY4k@X8d1I5^>HccUn:CeHUmC9hfd9HiV^TKA_1f?8GgO8majUP
ZVdLL@_n__caMACl6n@\QHEDe>HncF:bJeHXmC9hfd9H3Gc6_VKSf?8GgO60F^DL
@WdYL@_nPWWgFOY4JII0QH^;HVnmENEBqbdYhkdW5oohDOke0B>B\U8dnbBLdO8j
LC@Qb1cI3pT[Gi]4JJY^Q?aLAbMaNo<b=@FiZ`DB=II\mQQ=nj9YfUE=ZMN7]k5a
n3jno;CF\N=@[kD>K;@o>JdBARMaNo<F68FiZ`DnoKS>o<Ej[39G;0RRPiJaGP2a
nWjno;CF\NAlUZY5C@@o>Jdm2Wj`Nd>b=@FiZ`DB=II\mQ@`[>MbV6V20`EAhkq^
?c2A@\Bl4^D0T<j]mhP@FVjf^3X>l8;3lB::l0e53L^J`c8?YUO415S6DTN1\O[m
GS=[R7S@\e1Ik<j]mhPEhL_2^3X>lQEA4`G5]e5L`;47NNm@SE@415S6DTN1\O[m
\_ghk\EL\eAIkL9NM\[@FVj2^3X>l8;3lB:3d=EQ@GLG^j>JeBPqOUaBgGHYd]7l
`3L_K2oPX<:UQGodH0dK7hU6`6UCbH3OAZRjG^LV;Lg<YO^R@081XZFNK^Smim\o
D3L_K2MJX<:U_Go`H0dK7hR;O8G7iKA=K4OcG^LV;Lg<YO^R@081XZFN_DH;d1\g
D3j5C4o3X<:U_Go`H0dK7hU6;;KA4M;[=BRmf]4TqNCa7?`_k`NbIjd4begl:jdB
AN8LiknagQ>6T\NSBQL;h]l`V]N<_<RgKd0RKD]mWl?BKW?3@=JGhjdObgDlXjdB
AN8LiknagQ>6T\NSBQL;h]l`V]N<_<RgKd0RKD]mWl?BKWJ_a`l9fjd[73gl@jdB
AN8LiknagQ>6TKkXD4Og:2K5QBNfGqSQd_:9Zm7_jIRR\SZYOS0mG\`I<P;P4OTX
RF]8mbjB5`jBRHlHHKQV6Ejn\3jK0UR<hFa<6abgcT?27@E>>]7mGZ^SLNVI:7]Q
\j0Bo@<Hkf5I^8i<fWfQegOjMgQi9L6\[Ck1Z07_b\?27@E>>]7mGZ^SLNVI:7]Q
\j0Bo@<HjfoI[E1UH0mQeXOjMgQi9L6\[Ck1RnV@<36?:@ljV>2CAqdWN>6H_Ci[
YQBjkS970>k;LGJee]cN0LP?h;e^O_1O`6\?I3RFfH9gQhQiImoWFm79D9lMFaC[
]JJo`mb70>kC7E=Z7`<YRkD?fm[YAGGGV^E]X^0RiFcnhAmnbPe17nLiCH:P_oi[
=`bSR<b70>kC7E=Z7`<YRkD1X4ALAGG<`McWa@^OIMRnhAmnbPe17nLiCH:PI3l_
]ZWD72`1=o9R]pkK_c0LQ8ZTU:<I:fT]>05U0me>D34V<?\GVi`0nPh]L`acUW:N
A2A6L:@K3a8:9D@1VCNd=]CPLAbdJiT]F@LQjYGXJ6i4iSYjWgD>TPh_hd]8B3bg
;Gh6W7i8B`ok2bmOH2E\QjZiPAQ>0OUk>XNWjNGXJ6i4iSYT134i=2V?8LR5OSlS
8Mmo<]i8B`ok2bmOH2E\702D?@;noO@IdlKdXq0malokaUeY3>n3C>LLB1`b>TNC
`_B[V^XbmR1Xk5:Nf@maLQQdd^70]IRef>do`B<4ehAbSJ8I7807=j5WWO^SKo>U
Xj@ATYTBJPFFYg<4761^@DPBk:\XDFYM`^bc[0GN3UMoa0\QZH>7X6O>iQf@>d6C
>_aO\UaBj\mXk5:Nf@mdj\QBL5_f@]U2lT\4P_<4ehAbSJ8G7Y07=j5=I5^SKo>U
Xj@ATYT=VgFFYg>@56jjJ1B3\bHkajYMdjV\QM[CnngQgE3_hq<[XI3o\Pk@i5L?
A4>c4lTJPVmC@8@`CSiT?`387JERQTQnojiPT>TSXGCFWXjMCHlcfemgnghH6=eU
m2\>ZH@:W0Yl>50JS4T2Qj0fBkRhkic9Jg;_Lb^SYGjN[X0LAm_H<C0Mkf=dk1`;
gO:iW`TJ>MBDio11Lb5?i0387JERQTQSi^<LM7755?e4FJ;39@SWd`0;\CkA1f6X
TMolNXJ3n8El>l0JS4TlmP<g@]W0=lOc]Tg\1?\DKY8>qYZM4E3HOl2<ABmOSO6d
\HXfE=5fZAK00R[o?mf[PY=RV5^lf1a?c6__R=J1qFDGEQlbb_g9AGh6G:BC^8mf
U?JK<T1WA_FBMgieA5A1>QnNDQXONBDb3[J0hkFi>kDVNQOoKn]7;`4QLCf3^_e\
E^gRgj_R0ciJjiRI`5EX6JB91J7f<Qn6GBNn7h_oc?XFP66P;X]7ZoPm:ajD4ShQ
H77^5?RP[d8>dgieA5A1>QnNDQ5Of3eFL8C[ZSB2Jk;UK2XbH_JoE_olaY33e<gf
DXgRgj_R0c1X:klkVISOZkaB=7K:aQ:4W0RpFFKRd^MNb<D04m^TlkUUb6DjbPNb
XcQJN<2CFN9nZo;:i?i9Wghk^@7aeZ@ZRi?Di_;NBH@<DR>T:Z8Wl`QcBWRhL:HG
aco=62SkGXI3jk@m\6e2JJ71HSWXRiXLmLlBBHJ9<?naQ@^gLHYW@4PRD@Hd8^PG
hPDG`2JVFN9nZo;:i?i9WghklDQ67M^TS34SFl=BKmMMb\NNV?>GlX3O568N=:Hi
aco=6@RUSSlc;aV7mCI8MT6[f_c[i4q^26mMHBa^;M<XjZASL\B^RmoHEcPI<6Lh
d62RGTUc^EleDN8Llok2FF?[UNcfWZR:HEP4loPcHJ\]?lKd2O:mJbbmEaXgLiVn
M23Q?;LoT0]c1jm^mMeW`g5BMQ<k@KbF68;UMPCjj\XJB<?30n``I:5MV?nIf>BC
2<F6GTHc^EleDN8Llok2]Gm]S^>Bf>W[kEOi<2?^2O[1WOYSLVB2f:\cEa8gLiVn
FHFeLIndWU_h4X=M^:nOZN^Wmp;9i_7iJo41[b:7CZl9ZG`jUF;I<G<>_6M3k6Je
m<m1Hc;;H1WZlL]FmjZURT5HG43f1[L7JH8Y7[]ocAH9ZGaa6DoM;E<ZCGQ8U??O
1T8D29JIQ:`kWUH602F5<j\bdWZIOPNn9<2F<k]<eZH=VOP5K0[3BlF7PX5i?JS=
R@m1Hc;;H1WZlL]=[[BDMJ[;mCT1D5`m=3BXbc4\DAlEXhUgKJoM;E<ZCGQ8]?lH
5n3RQMIR8ebc?bbg[RMQpd:jDbASj;N4Fl02LSKIXXZZW991kXY2lD@ag@iKEach
AZahXjHllaLM04`aoBPe<Va?fHE`_YVHkmFiORKIXXZ=Wo?;nSEoQXV9jh4WTi2H
Cb<a`cHg6`GZnG<aETUFMIVj4@>EUVWVdeY:io8AjJY>SQP^=7_:30amCHl_6_ch
AZahXjHllaHeG77@c4S1QY0djGX`l7O]JNFi4Sc>Kn6^1o?;nSEoQXV9jhl4D5]G
^YA<K[LC=TQmRo0p`;lYI4SHdXX`\OLR40:b@[f\PL6Df5UM]=l3]1gLJ6o9hH4>
Xj=TVX\=QPd1o2V7f054^@H6CTP4f7_RW0:6@[f\_CEXXFgUfC_g3XZWmXLi3e?n
>j6^GR:4@Y;@\VAf?_\dnbR`F;V1HZON=oNcYTSf@c?3R`A5?7i]RDF9m6kIgU4>
Xj=TVVN\M<NY0@E>Hk59B?V\dXITI7_2W14WebNB_CEXXFgUfC_g3XZW;E3O7iFY
<CV_bMTPE_q^V?daiN^KIo=n1U>3JIOF^[5K:f@h6g^MQDU\mK>VFToPU?3d7`hc
Ma9k6_;YXQ5EDR_E^Chgj[E31U>37KU_8Z?2mH7c6`;W@IHGAO2>1MallRAo6S4U
lXoDlDXYdQkD^@IRVJGnLBcneUAQddSNG\e9GJZ_3?NlbX>\mK>VFToP0ZPkRN?_
Ma9k6_;8Y_LcMDm?>1n8b<H<fSVNc=Uh=FpPITgGYIJ>DUf9`UCa?8kQ?lUh4eE>
f:c@^nq]^aI9hhfneLnQgL0]`<9h]@7J8]k=BU5BK[CSiU5^g<WY:LG[:JWlWM5e
I?0Di5P]?\I63kbHN6fdZSKL@^YlUR[WHcLDjU^cH;K]?YjO5maeQnbhX`SKVT[e
_eo>V6O_X[\bGcG[U6`dgIQg0Sl^D6aN9U3_9MB`AaQSiU5^g<WYYaG6h`@loBZP
A`=2<gL8ga7QFEi@gAUg5:?c;:CT7Uq>1N@mdZ\W4fd7DLl19mXQHlEELIF34VO?
^G@Z;Bem3n^k\GG36EDdPe93BNMYXJ9XG_TUBZ9W4fd7LkDjiXQNdllfH_D\2iS?
d:23L^n1NYDEk2=\RVAVXgDOh0XBPY_;iZeY\^644N7W<S0F`4g<=^`OgBmDh_6[
dG=Z;Bem3iOb;4c3k`PZ\BZJCI7QMLj1G_bUBa9:B4JTI0jB\]^5Reqmc8OG]McF
AT<jL0FIWWVia1D1GJ@=FBR8>@e;;YU7b159nI^P75bE`ed=382Q=:`PUGg0FMNF
AT<jL3:Jh<=i51F1O<dZXNa8>@eh?>4_95V[M]KacBl[kkBfBfG9CDK?X9Z<LS38
?Cbb2W;FljCD?3^1bg8h_[J8>@e;c7XV\\c=nI^PhSP2LU8H]B7Q=:`PUGg0F2@3
_djI>N?0jkA_Y5pB_3Ym_A[?IZZ5AJha]hNe3`4W>2V2VH@1MPKUcK@U3V;]`KMd
b2l1njeReGhUfB>VYQ9jgAf?IZZ5AJh1af5^kCB:V6Q_[Vo1MPKg<IBCm0=9bgfF
PaYS2I;eV0[I>Pa3?dchnoZ3n?IGRSX_ekaDfAN]8<bXVHd1MPKg<HBDoNk]`b0F
b2]1njeReGhUfB>VYQ9jgmfW[aBcOcDmIdjhWbq7]S:?Q]C6bB[K_VnX0iKdhnE5
aTLG9\CLa_T\BilMRQZT2UTVJm8f7o^`5c=\n1]ehD>@e]`6bB[K_VnX0FnJ>nNT
eLO5R\@IB`Qm;RIeXQbT2UTVJm8f7o^`5c=\n1]ehD>@eOo1H?CNNVdX0PnT1\Z@
4`ZG9\CIB`Q[@Gm>bYA2Z:LhUkfq;4m;oXH>fR_ThlXGqhE1EmTBj17\RgDNC0eF
aNhWRDRY]^YNN_8^O?<`6[^P3GQljM:3@`MHl2SEWGcWnORU9V2B31WX6Se2Lc>\
GGfW@DRQHPL2I;1Z56oXl[^P3GQljM:3@`MHl2SEWGcWnORU9=]KO3TbC]DNC0eF
aVl?P9ZM7?L2I;1Z51@`WhKK?3E\=09BmqBNKM2hWc=Y4DM]2G@F86Yj^GM:PE?[
>BnUbI8RWT[_WnRoO=FLYgI`8`QEYmKgZF@ED24e9\Q@Jk@Y]Q=QQd\V?o<McE7Y
j4Ui_XoY19_^YeI<j3Bc0i<n662;]ET@6U@ED2;HWA=Y4DM]2G@F86Yjd=lEkU[h
SX0EQ;FOTg@E_21oO\FLYgI`8`QEYmKgZF@ED2;HIA@_`3B[E@]0BZ1^9qOUaBgG
HYd]7l`FoCC4o3X<:U_G80LVl;\7fl`AUfbH3OAZRjG^LV;Lg<YO^R@081XS8P;^
SmiW`dM7IO6:260dGAgTl?Y=<4chR37_?BP59K=Ibi8Pk58D`7QLB<dl;TXZFN_D
H;d]7l`FoCC4o3X<:U_Go`H0dK7hDR?c?XTQ3@AZRjG^LV;Lg<YO^R@081XZFN_D
=h;DB:XD;c6d0`PjPpTP>[^L:3C;3@hd@=8IjCIRN<PG5]JeGX?WF6Q73J82RP3H
h0f<R\D]4e6T=>_;N1=g\]^4O`4Fh6dYnVQ?gKmW:0N]FcDG9896noIP9>CUPS7o
m8BJjZ8M4aDB8IYOg0k9fk4N:^C;3@hd@=8IjCIRN<PG5]JGVajWF6QPj`C2R8nh
8:S3RbD]4e6T=>_;N1=9f]4NE\6MS;Vfe2j33gTMhq0\g6PFUKB65HSbN?X:gJ5F
[U\F5KFH[jO:8bng_KL_LnHiij?VHT3MJ3YLEU\IC>9UT<f]nQ5DWIECUjN6d=>8
L4Z>CXO?M>]:jnkcI1I<O2dkaK_fQ=?W6j6c;0C<Lmn9MEa<UUB65HSbN?X:gJ5F
[U\FC0nlFgPFARng_K7ONU36oWESW:ERH6YLEU\IC>99MOa<R5KnNYm?AWHkfj7_
Uqlfdl1[gLW81iePB0B9TGA`]JDR;X>SRM<;dVVX9hHCkZ@D8J0F]IiOhQ>mq@J1
dZ3aeGDFCDEXCTfc\TLan06dMDB=;X<iZ52?Z4d>0oFVD4JMVU@IW8_G=WBgh7;R
UocEQ1=S:i\NIlmEkVA]IkEKYDB=;X<iZ@Yb2hd2liMJXh7i0I8FE__gA@5UY:i=
8m`]`7A@ZVVGAlKED7635C3ai99PKdX>jNjCR3\CkJW7P;VUaG5JW;l7Yh<`7@dF
LFoH;aWFCDEXCTfc\TLan06dMDB=;X<iZ@jC93WIB_IXGfmQC^=li51qD?QMF?TY
6;0<EM]QAShd1:8YWT3XMQ[K?5jMj]5h9GKS@AK@NIk`=k_Zf<`Q<`0SUO^8mMnD
>WQbU5Z2Uk>b`Yb>fl5@@R[S?5jMjZbWT00QIjcf`_ke=NO7b[o?d:_TR>1ICeg2
6NQPUQ[7n71K1:8YWKg<UB56[o_>hdWLP8><oI?hFI8JTAGP2[GG<UDkfW2RI7iC
C:36ih4;S@DSnd<3fl5@1FPZJ?kYfnP4T0cQO[`ZL[hjj[6V7KWbRP^VJbCZYhT]
6;0<WjL3b98A=C>NJFKeq`H\G`O5Q0faWZJ>B9;n`Y4FTJ?h8oRmgeOYWi5fQITb
jHOSYL2oF2J4`C@OPej:eL9`OXc11^j9S;Q0h[[W>c5K]Ig_R3VmHeOYWicWeZSQ
dkWHF6NgJY=;8@@R64GXTEFGOGP22_Fj9InmAP[B>Y4FTJ?hcM`UNfN[loPKMOV3
?Z:?mLGo?2J4`C@OPej:eLW<7E4SkGFIUnMkBnJfeL`gYjRC4HneiPVC6X>31ZS:
XXSeoLPfCVU[[FEmKEL`1K5]JfD5J0faWc3=aGTZO[c6H5_BbqL0TI5B>hmcP0Ul
62ncOmfl]4IIN>:lH`2H5CY=\Qn]Gn0IYfW5`c6aVV?ch5_;PVfTjcX0jUK\4:8K
:>WI<d5N1i>;M>ONe`J8h]PZV=o_oUa;o`7_gh^SKojh`X^P5akC::LgXDZ^LUBC
fQ^Q<dDl]eII00`jjZXCTk9oG?3>g^?lSPJ\UjZPV]4hg=@;39m`k^GA;@k@jE2K
;F40l^5l]eIIN>ENDEV\TbHBVoo`TioDgo[3bl?iT<0C_^dR]\Y8H6c6>hmcP0=k
BA;8KgfaXGHK;DpYF1;?]YmacAaQ>:C4QYjKdOYHFg:\J6AWAbbp9Fchc`V<PG5?
YeT69`E=a:>9iT1PUGD6CDEIdTf3HTLI]kE[bLe6NH08]`8oG80NWYajo7FC8D9E
Q_F=MCYGKI;CmlOnZaMNO7N\Z[XO@>;911=?c9CaNl0PJO\LPYC[a\fEWIl=NIMg
T^BB@WnWC4;om>mIM1=46e`^QYfjHTL^_Z3Cc9\d:eHc`Q8E>YoBlgMC0\hEnU@N
P_ACMo<G]@dgVFofZaMNO7N\Z[XOYnA?:kE:bS6_6dXi0Oj3f3\[aJW]^;VhPG5?
YeT69`E=a:>9iT1PUe18HmYfo?dFW6XVF^q47Z0Zl0Pe8A[9K;lECUi1]EK3oBOV
h]8E_3:Ofcmd27Igb`>h^dkI6A7b\56DlVl46c_7:R^\BEWYe<AGjcYc;]N2Fd1A
go5<\bm<aBTe\_F`5X@L^ZEXSMMHXo1Qd2]hA9h`MdhaH=<NoE851h12;c<\5N4g
AEmA^cjmn1bc`T\1ToP?DPP4gUih=lhCT]h46c_:TRNe8A[9K;lECUi1]EK3oBOV
h]8E_3:Ofcmd2\Mm66`Gnl4heDELjmqY8QV[3bd\dk=Y9D5hNK@:h@Vb5GiZG>17
T_IEkUgBnfWXbY;O14jUcFBZ@0K9<cNATD8k]6@m_Cm2QMg_RV@g;bRC5KhF9T[R
FcNahP@XJDd`^<LP]ZgOl@:f_4U4P;dU?6_O;le^GC8J_6BSl]k<VcP`d\@Ue6SE
`SZeHmiN:bF>C9nO1MTLMOB\=LOm3g8ki8Rd7bK\dk=Y9D5hNK@:h@Vb5GiZG>17
T_IEkUgBWV;EN<nkc>CnMe4H3pBj?GZMkgD6cle\Z;_fVKfW;1OHL?=hC8hJ0:6G
>C9AoU0d]k]ic^klI[QcYm\hNAPP@_DXfOeOJ=l]]GXO;EWf?ZhGcO?aH^\cjS@9
E4mF`2VSbhmN5jE^JoU84m9n2mcSldIiDYo:O]lk[H0;=TF30ebHgZ1L]AKY>N6l
:FiaC7e>98]ic^K?odi8=24S<DiIYJOmkND6cle\Z;_fVKfW;1OHL?=hC8hJ0:6G
>C9n[fSlkA2F5l2Z<\^1pAnP^?cJ[;]_Pbl:R<COZo1Z<@Q4[Nm;gXSNVf^E1=LP
X7[H8a;3aGOQU5]VIZI>9^b3CM;VQ^RNX<;`24AHHXX68R7??iVY9CegKNOmicLo
BoF6W9:7I[N@f<_l=33eK^a1^o<Y\HQIbh;<BVJe^Tl5oCS5h?UkZblUf82lZoF?
T6\aZi;3aG`kG;@a1=;>ZU8[k>lJ`;]_Pbl:R<COZo1Z<@Q4[Nm;gXSNVf^E1=_V
M;QBgRRB?>FY`=4pK5iP??>O9AoU0dbkPaLT6^JmU8MNhn?RiIYJOmkND6cle\Z;
_a@XZRXB9CHjb2G;DKa9?5<m<nB0el59BC]h8T:\e?]E_e46_k7J1=DN_:@GWmQJ
0;llkW;EOHL?FSll86RiLONg9]Te?l59BWcmR5`?1HUgXk9ePUE:[4_TVlf=FR;M
gVQ9=f;`OHL?=hC8hJ0:6G>C9AoU0dbkPaLT6^JmU8MNhn?RiIYJOmkND42e`C49
2ZmR8=39c2q9`j@ABFLT\\S0kjlA;5XG^81`S5Q2BghF5PCYVbV<Sk94^iGGeQHJ
e]FkE9YDR^daDZnF?>aML]>2Y_A>7fm^5_EWPe>d[bCfFa=93^c]6@Hf^9;;6Z]X
>7kP0>Q3n:A`LX4c?3fZZ0heY_O>W?U8ckI`hAY@lA>?n5F_LFElZkm4^iGGB0@6
>7kP0>Q5j5AKG`=mUF;T\\S0kjlA;5XG^81`S5Q2BghF5PCYVbV<9SH[omOMGD9A
m3<Qjq`EMWTeGOV0bCQjEk:FaZlhN@KKNBW`cg]CFE^`e22engI>2M]13fka=`o3
R[giA61SbZXDCLL6ZH[==:Lad\O:OPi]I0]4=6\RhFneNn\b\3eF2PoG<HElf<4l
Mg2BSWkX4><0Cmc;d]MY=OLaWLU2GEIKBC<XGBol<I5TH_cK3ZI>2M]gKVGVfH4l
Mg2Y_fSkQkK<GiV0bCQjEk:FaZlhN@KKNBW`cg]CFE^`e22TOmT0eE>P3=`QS;L]
qP`6Z=h8]5FTGe_B;i=Bjd;d;pc=[^ck9Uflib8bnR6cM:SEnccK6LZUHW7`FAP;
g=c82Y4IdPN[HK>mOSf;2aRNPJ<lXnjih4NI:;i:FGFi\8`H><UTB`VaKYO1d<6N
cgh5aZ^4=hSnN1L4R\QD8Rd92g<lHE75=j29e7H:FGFiP8L61cJ1?448DI_[3lSU
iBn]@^4IdPN[WHj_AjQD8R@FX:@DFf];9Aflib8bnR6cM:SEnccK6LZUHW7`FAP;
g=ccif5fB4^S3F<NBoe2pU=5QbD7encMCkk6Gi8YdIcMFK?>eQKIm22NW8^oJnF^
0EK:@OhC?Eg_aSVfU_>14Hd:L38of6Vb7h:<KCYkom`fh8OiWH6c7<k`FGHdDf<C
HZiHYRffk=ebA;GAch84DEdN9kkR`ecM[kk6Gi8YdIcMFK?>eQKIm22NW8^oJnF^
0EK:@Oh6YgMQcI\m[5VFl4PU9Qdm:N7<3EEjOogaJ3HgqWf>jJ17B;0CdM]klShF
k:8jST3J8Q[H<5jJ6]5f3GaRK[`k?[hk7FMCliZJPU02O5P0PE_fQ0GM9Kl?@cQN
Le?^\Jaj^RQL^P0P^ZAgcVB0UgB\Ac_^]O_:oJad2`h4LQlmQ7i\4>0C2M]klShF
k:8jST3J8Q[H<5jJ6]5f3GaRK[`k?[hk7[6<kKWUXP^VbbC_@hTB=_nc2^4^?g;T
MFlfp<SHfbJg0Qcfb6dW3o^U=J=[<biEPK9G3a9pOgRdc\kA6Ii1;VNa@Lgn^`^Y
Af\O;@Y9ieDQnem56HX?5n_CF[[D_GfQSBWX`;@jBik>`9KDONB[nl`YJDl`kO`[
aQhmKJAK2OAaBfk]JfK[]ECGi[;90J<2SBZS5idfOTG2Vf9:@IiZ;VNa@Lgn^`^Y
Af\O;@Y9ieDQnem56HX?5n_CF[[D_`]TW9CWJ74O^5R:_>_9A81e3AKk71a@\9jq
O1;6EWOASQO=mJbbmEaXgLiVnFHFeLIndKY>A827D21g1`g6BMQ<k@7[^BH=V=o3
cH>6eXH[3YTc79ZYcmkbnQ[0>doeX[1h6Ae9Mb2WQmMeWE\5Y`76?ZQA^BU_R42K
^2O[1WOYSQO=mJbbmEaXgLiVnFHFeLIndKY>A827D21g1`g6BMQ<k@KbF==kiVBc
^2O[1W:Y@K=KJefJM7e955TqVPPVZa?ek@4PbHcJ>j2Q?m@PlOe<B^Wa?>_9\]ZI
Y33=6l[e[CP\VQL:Qo9\FQZQ5gJdf`kEMihNQnIDoZioP6?HEIkgXDXGPdgjikdS
NKGNO2C5X=KM;9LT4J8lTj4IWbD@Z@?Ck@4PbHcJ>j2Q?m@PlOe<B^Wa?>_9\]ZI
Y33=6l[e[CP\VQc:4J8lTj4IWbD@Z@4ke]leWHfgIE\iP53pPBf;4aLCXZ893T5V
``U;C>]4IUNSN;?LVAJ<4]ebXSYFXIHl7_E]0:jbbcTjNFIRPOGmiF3DgINWBe5F
``U;C>]4IUNSN;?LVAJ<4]ebXSYFXIHl7_E]0:jb[f_RCEo`Fg=AC_LCXZ893T5V
``U;C>]4IUNSN;?LVAJ<gRBfHaF9foU5@gVlq=D4j:KE_4mY8RY\_eP9h18afSFB
70CSASNXkXg52YL\k^IF7MoO29W94Q67I8<NV4mE6kDE<4mY8RY\_eP9h18afSFB
70CSASNXkXg52YL\k^IF7MoO29W94Q8c<o33J4mE6kDE<4mY8RY\_eP9h18afSFB
70CSASNXkN__>^RN;>keRZeENq4YUY__i@VD>:8l;gKHT5m1_mjQlV`MhlJ?9m\3
l778diMR?Ymhc@Lh7Ll9Ya:`=W;_3U5^i]VD>:8l;gKHT5m1_mjQlV`MhlJ?9m\3
l778diMR?Ymhc@Lh7Ll9Ya:`=W;_3U5^i]VD>:8l;gKHT5m1_mjQlV`MhlJ?9mSO
@;\=HJ]h]J3OYeq>_kj8n2]F@d3ME[8V9DJ7X2\CUh:2:S\?[n`KiRio>N`BI;dd
kH5fD2?6U1]AYcODMcGlU2YF@d3ME[8V9DJ7X2\CUh:2:S\?[n`KiRio>N`BI;dd
kH5fD2?6U1]AYcODMcGlU2YF@d3ME[8V9DJ7X2\CUh:2:S\?[n`[KJG_kULjN7i[
F<=S`q^\Q@g@[DPo6O23L6HEg5@b5UQb4]kk\8_7a70_`2haXn53\h\[fM5U8TgX
QX`Zcj=EE6YW=lQo6E23L6HEg5@bCnmUFPOh\<_7a70_`2haXn53\h\[fM\1_<@[
Taki4W^6_hG9[TPo6Oe`L3g<jmQ:YM`SkfMkqdBikHAn];RCaLN@cK4THRb`eRJp
Uf<Tn2\?:]ef2PL7Q;=B?akHSHU8=h?cYWIS>EKl4[[bO:KS7b4Zf2E3TImgcV<:
nkoL4[\l[>7_UPHWH0=Q?aU:?[n[5i?dYWIS>EKl4[[bT5<=5DY6_ab]T8MDXV0[
U<;7=:\W:]efiOLmJcUUodkl2kEJXep6FRi1UO<8m\h8egCBo=2FXC^U^nb0ZgYS
S^aIRUDR9MAL\<^SI9Ll8ZccUSfigZ8KA0MK4kihU0KU954P1e`GmYZA>dJ<QLlQ
aPjJ<XfKIMU=R3YWI95l8ZccU7fUm`n6m0:K4kihU0KU9Q4n1PZJm^NA7C=Kc;>4
LP625QW7h2U>\cl7?0FKPCTL>YDp67mYR\J80C0LXN2`ZHlNSA5@enhT`[CRo4l=
IJLOfPEbX9:3QLL^IOX:\OecemP1cTn[lYJ@0C0LXN2`ZHlNSA5@enhT`[CRo4l=
IJLOfPEbX9:3QLL^IOX:\OecemP1cTn[lYJ@0C0LXN2`ZHlNSA5@enhT`[CRo4l=
fEY3g];ToeFJ8F:bHmqQ5\C`6B2AJIgN61h`op<TVhY1_QJ6qL=;55Yq\C4R94cB
>nH7lHhY=6pgPnTU3L3=hC8hJ0:6G>C9AoU0dbkPaLT6^JmU8MNhn?RiIYJOmkND
6cle\Z;_fVKfW;1OHL?=hC8hJ0:6G>C9AoU0dbkPaLT6^JmU8MNhn?RiIYJOmkND
6cle\Z;_fVKfW;1OHL?=hC8hJ0:6G>C9AoU0dbkPaLT6^JmU8MNhn?RiIYJOmkND
6cle\Z;_fVKf^@eXTSLdIYgkIR`R<qmScQoVmJQ^DQ`LE=Mfj8<2@PkVNFGmd@c7
P0F<b5^XRjWRC4GSRe?EGBIm\>B48[RB?6pIYPFS;Idga<E`<mbaP]\kFKYW>UgT
G01I]EOLePZM2FLH3?`hP8TBO3GMGHnnB]id<\1oGIPga<E`<mbaP]\kFKYW>UgT
G01I]EOLePZM2ch9T=AG?J1=QXO_GDRnB]id<\1oGIPga<E`<mbaP]\kFKYW>UgT
G01I]EOLePZM2FLH3?`hP8TBO3GMGHnnB]id;c3ef<f[PDHV\@]S1pIlHYPnabiU
PH>eM;aB;]VhVSWjKF^O;4k_XA4aZ>8MPcHmLl:mWOJ^6eGFE\IRB5DO\4?BeM:6
^To0Zh8B;5VhVSWjKF^O;4kgcC1:KH6XeabjS71QlRf`3LGA40lQB?h:3FH_aciU
PH>eM;aB;]VhVSWjKF^O;4k_XA4aZ>8MPcHmLl:mWOJ^6eGFSP7JcohSk3_UeUPc
:@Z;2;VnpZ09T@MC3EQNZRNh[U9iBMDKeRQSj5<>Be2KD0YjTd8gmQ?nP\6T>>[A
<<7C:lVI0ZdQ]oGGNh[G_GPDcUPbY6d>S[0LE5<m@ISA:K`\LIBg0Q?nP\6T>>ki
IjOTCPVIgZJ\T>[C3EQNZRNh[U9iBMDKeRQSj5<>Be2KD0YjTd8gmQ?nP\6T>>ki
IjOC35G?c]RAWZYeklEYkCUYAR?q^<nbPMOMUDlnfZ0YI5Xa>B=B1oiXSknDQ5S?
lYAUMQ\?\oD[7kI[]8gTOaokMB6<bn]ml_OHUDlnfZ0YI5_F=LnfAP^lcKEbN5S?
lYAUMQ\?\oD[7E>NP]UhnFk<MBYle9JY=>OOUDlnfZ0YI5Xa>B=B1oiXSknDQ5S?
lYAUMQ\?\oD[7E>NP]UhnFk<MB6<bga<^_YC<jb3edoRZlp8\n>Y^RQWFLUPQQ@e
520ZXS3hoD45i5>deEdi<VFBSejS:FRM=bCZMXYT6m:mMLimWYj:2RQWFLUPQQ@e
520ZXS3hoD45i5>deEdi<VFBSejSXd6@>Edb8XZT6m:mMLimWFj6A3cWFLUPQQ@e
520ZXS3hoD45i5>deEdi<VFBSejSXd6@>Edb8XZT6m:mMLim4jm;RB@TU7\^f21X
KqX3Q@GQh[^V_mTm3_eVXDIokQN;VODd^^7ib0R?2E>hGK2Q=Xk39WnNASnj3>gb
77blLn]DhG^V_mTm3_eVXDIokQN;VODd^^7ib0R?2E>`Feh3m@:993nNASnj3>gb
77blLnUZLEfV_mTm3_eVXDIokQN;VODd^^7ib0R?2E>`Feh3m@:993nNASnj3>gb
77b<On?aZ87O:f63j:]Pqb419=XA`LDHNljV4\dTijjSLU]T?OWM5N3nOVRTe[ol
L=MVD;j[I<4M]l4FGV1^gKR2j11AYLDHNljV4OZTlcjCSU]T?OWWFdg@>VCQ0HSX
f?WN\;J[I<4M]l4FGV1^gKR2jD`OX5DHnljV4\dTijjSLU]T?OWM5NTWIZ`Q0HSX
f?WN\;j[I<4M]l4FGV1^gKm2eEL2Bd76k1X5IaBqIQc6:Z<j_\Snf9SXZhFlQcgm
oV[6^CLbbX7F<P17_8D?<Zd`Ro?6lmeUYM3aYJ\:IDm]nk<h_\SnG9m]ikK@KcR2
o7i=i9LEb4H?<A>;c`iA<aH4`P2hQBn_YM3aYJ\:I2nTg[8TbSSVf9SXZhFlQcgm
o7i=4]><5X7hTiX:<`iL<Zd`Ro?6lmeUYM3aYJ\:IYKZDjj:T@O8hOYP>nqWMS0P
4CE@d4@eH`LacG4k8:Mf^M9m]lbnYH6eTiSKX4ZI8nQJf[FnNA@dV95heV;W9ecm
2C?@d7APbdXacG4_Dn;XY>IQa\kA?HIbCTg;C4ZI8F4jf[TL=kELVT<nObOKO\Ok
\IOG84ReH`LacG4eU<_XY>I`@`RU?HTeTiSKX4ZI8nQJf[FnNA@dVTlnObOK_fYR
LBhS8V26aQU`?p\jcbX4]U^I9^Q0lioo]nE;T[ZPb74FO;3X8PF0c9AJThef_VQ2
1@ifN1o`:2L4SM6PUjR>`pXSDPESWjdDniG5;]A1YjBNaCR8Xk7KXG46FJ=Z6RfC
67eCQa?R9i1AGnjj>IfU8lLR`=QQ^jdDei>mHX2GTUQNoRF8Xdh[I8D6FJ]AWA3N
6WnMlJ]0iCTA\5Yjel<AUA`COk;Cil@]nDG5;]Af?4`X5>C8Xk7KXG46FJ=Z6RfC
67eCQa?R7iBD8XjjeI<AUA`f`4VG_9>PDe@j33:Wp?Y^gnXYg?LCTld4VEon;Ie:
M02?KKgSAj50HmM;X]83YnS3ZAjR6cM<YZo`5MlR5Uld:N7\T>LCclmXZmoiee]X
2g2?KAIBg0501bAIV_@KGn56N5=]FWRQVZoJgoC?_:7oLMfPECbCTlFGF_H=M6g:
d02?KKgSAj50HmM;X]8?QDIM7A=]XWRQVZoJgoC?_:X2>;UTMUDRD1SeoSTq<mB?
7h521lYRlENHijoif7EBBP]<4nFk_MBGKbn@cl>gkh3odGB\oYTWC>Bed\OH<V[j
L;c`_lYREWNRi8oHKGb87P]nHGNB`l93e^9XLlaZ]h;@GfZfGf5<C>BeD1og2Skc
MN<0W3Y<@MQ^b\oOf7EBBP]<4nFk_MBGKbn@cl_WmUDG=fZfZI5NC>BeD1og2Y0m
[FYC?TS<e]eSYQq_S7lbNM[QeH0i]ioDd=?]W[<D_Clmi_GYUGFHSZ^KC[HC=`_6
>@SRk]Y613<2Id1_e1iIN1lhUYRi]ioB5=3j_<:G_C^miJbXTeRB:ZCKC[HHUF?A
>@dR?ES613<2I\d<6hgI;lZhPYWGB\l6d=?]W[<D_Clmi_GYUGFHSZ^KC[HC=TAR
YQ^l>\M613<2I\d<:j>nGDK:eh@;:UORDq8Fm?]I]4eFj^QG[XGh;O`ZiMP]kIIj
gG=:5J_mqhX;6mhX`W8`PVQmaN;WSj3QHfMcAAEBcg5P\_l1@oRk<nFJgJkhU\mi
IcKLkIDDVh878_8Eg?8Pb<9:iG;W:j3QHfMcAAEBcg5P\_l1@oRk<nFJgJ5OVg0:
OcKLkI2CL<5BF[S?m[EPS<9:iG;W:j3QHfMcAAEBcg5P\_l1@oRk<nFJgJ5aVg0:
OcKLkI2CL<>0ZRhe;g[7FY@2kVIpBEohhXP:^WNZaiBSi>ik]\Go0N3NG\_>6N:D
Ti`NIY9VQWNRPlO51e<4oj\F<QSU=JOk]jP6^9HWR9Zbi>ik]\Go0N3NG\_>6N:D
Ti`NIY9VQWNRPlm=d[95Nj\N<cKbTE472AEO^9HWR9Zbi>ik]\Go0N3NG\_>6N:D
Ti`NIY9VQWNRPlm=d[95Nj\N<cKbTfdaCk`hdl`O[gM7OWpH3U1C]7Y]>TA<`7lR
3@`VPDjM6S3kgK374fN`kI;hhbj06M^S4BK4A>Zi8[a\]?;A6XV\57Ae_i1a`7lR
3H07PD2M6S3kgK374fN`kI;hhbjdBMWS4BK4_hJZ8[5\D07HLm6Qf7Ce_i1a`7lR
3@`VPDjM6S3kgK374fN`kI;hhbjdBMWS4BK4_hJZ8[5\]?;AK]BEJ;>W;:iNT^cU
Xp5j^iIX3TP=KFiVZ>a0iLN3L9VA[46:JBoJ<?@0`Hl?i4WRF><S0XMEAZ?e?bnW
38WHoaj[3\MU6hM2ce^goF\gMQT9CUg?XPIJ<;@0`Hl?0PefbHOS0PMEAZ?e2XTk
ja5W4\j[3\MU6hgVZ>a0iLN3L9VA[46:JBoJ<?@0`Hl?0PefbHOS0PMEAZ?e?bnW
38WM`GJQNYg70HVADk5npoeYRH;ocHBZ3d`i^@VXOV5`hZ?0F^1?lj[UihL58AMQ
TM5LDSFTA:;;`[:UB07^6lamEhl\o4Bcc7RCX7U90aoPbL\K2lDmb5hn^DVXGJm\
O\6RESFk7ZBE10BV@HXdKlamEhlo0HgIaR`i^@VXOV5`hZ?0F^1?lj[Uih4@>lMQ
THSefNFTK:;;`[:UB07^6lo7VfUh0elPi^RXMLPpmmMb5eeR3U99_j1?ODdCbMRT
oT6?IZEg23=^W>_lZ[?n_]N64<=H^WJ[8cb^e`BQ2Q7[ICmXZ0i]]j1`ODdCbMRT
oT6?IZEg2hhbD=M?Zj2ZagE1hPQcSXjcma<Ve`BQ2Q7[Tken<l2N]j1`ODdCbMRT
oT6?IZEg23=^mFe0db?C_]N64<=H^WJ[8cb^e`BQ2FT1Z2HEIeOUmH2;e1qo<DBS
:>SP5=LP]j;U2KAPMJA]nMJ@N1CPPZK<[:Zk_ca7fK5cK4;G8jAgiRo9ANnT]IP6
\lHPZ0X]]jaU2KAPMJA]nMJ@N7^j\C]<[:Zk_ca7fK5cK4;G8jAgiRo9ANnV];`:
C>1UZ0N]]jaU2KAPMJA]nMJ@N7^j\C]<[:Zk_ca7fK5cK4;G8jAgiRo9ANnV6lNC
[:AmDbFEoKBEJpF4SioOQ\<7`6>7jn7MUPWcAMIGL;O3HKo1IMOS:7aXif_=NAB>
RbLedd`d:?P=10Fe[P_oQOjGH:A7jY7MUPWcAMIGL;O3mUaS2POS:7aXif_=NAB>
RbLedd`d:?eM;AneF<PoQJjGH:A7jY7MUPWcAMIGL;O3mUaS2POS:7aXif_=NAB>
RbLedd`d:?eM;AnB3Xa24jD]g?P7YbmeqkncH1MlUBGF[EWX\@Ck[<Z@RlZ\;CbD
I1a;l4o4Y9jfU:ngZh8a\4VbW04FmX4a0PmZIDBp@QB<7WTBY<mb]eSOUocZ66?F
ojFg2lTmJVg^\Z93<BW_26\V96KkM]hQHfGcf`h?@MMNGeDRbK4QjAS[UocZ66?F
ojFg2lTmJVg^\Z93<BW_2<lVj6nFHcT<f[mO`bGmEMfF\ZTJY_BZjAS[UocZ66?F
ojFg2lTmJVg^\Z93<BW_2<lVj6nFHcT<f[mO`bGmEI_`Ahd6d@28^AL6WMqZoV8A
G47;beL8G];BZW>=KibKIklI<b77\1YOZc?09fUMMLfO@ChWACMb8O0<>MZZMo4m
^Ek58eMOG];BZW>=KibKIklI<b77\1VGCPHmV[X0Q7AZZ<^F8YWI`\;i0e9Go7X6
I4f;bZL==]hBZW>=KibKIklI<b77\1VGCPHmV[X0Q7AZZ<^F8YWI`\;i0e9Gn>db
VJLI]VmSeR[YTqS74n1X[a_OY^SWCOJ74O^5R:_>k96W>^FP1B?WheBB`MAfCOSD
3UV>P8@AB=nlm`SJj54WE1:JYcSBGXJ74O^5R:_>k96Ii1;VNa@Lgn^`^YAf\O;@
Y9ieDQnem56HX?5n_CF[[D_`]TW9CWJ74O^5R:_>k96Ii1;VNa@Lgn^`^YAf\O;@
Y9ieDQnem56HX?5M2C^V]YJ1Om9lU?;hpMa>iKVQW`2>gl\XZohoRV5iaQVOc4bW
k\jS`fSXlE@>faHJYll:]KL:2W8AIa6m=MeJ<oET7ST>hlCZFShoRV5iaQdeBVi<
RZBS^fSXlE@>fTb8`?T6L`mMPJmW?X:24\WFicPQ6We5kEZX<ohoRV5iaQdeBVi<
RZBS^fSXlE@>fTb8`?T6L`mMPJmW?X:24\^A<9`T`>2EE`c]bRhpK;8QoCO1V:\S
VQO=mJbbmEaXgfGh26<PeLIndKY>A827`mMJWE\5Y`76?ZQA^BH=K\SEODMeXj\A
85nnBAbPmEaXg6X7>RHZeCgPmVKZ2gS`H]1A1`g6BMQ<k@KbF==kiVBc^2O[1WOY
SQO=mJbbmE@_o6me<RnIeLIndKY>A827D21g1`g6BMQ<k@KbF==ki@>oD_Bi78k5
g^7F`LqUFcTaHA\1lS[k^X8P7DVjf6L17e`4]706nmLm5Qk]>Vb1QX4hXV[nMH`7
ig0GFOOUYEcO?NhZl=A7hOSWGkYPL9OT7edDfFd6HgK>YLaG=Sm1QX4h=9MdmRT1
M4gjn28IYE9Q=A7O@==]^XjP_he^L9lT7edDfFd6H6P:oQh]3XF1Q^`lQfodMdf1
M4gjn28I_IHi14DLV0Uha_cN`pe4hdWI5N?i8C_B2CKARaXhI<PC\aTEdXcHGlL=
F`VKjk53Q1jj1OkOQ5[PoA\`m^eUH3C7\aAiV`e`fFh:kP6hoL9CE42d3[UVVBF;
VQZ[XJl\]Jjj1OkOQ5[PoAF6cKX56ZnE5;W`4<\B4?_:ki6hIRP9]R0eV1A1UIZh
fe_<iQnMbVQEaD_b6:g8YL`_3<XJ<l0ikRAM_I^e[mSmq_Va<BKe0_lOCkCL1l3^
:G^GY:S@hF4Tmad5>dbEM[e1F[FPL9G\7^:]a\IYZY90^_1EGYbBiflnfc`k@]c^
EdK>:[S@1F4Tmad5>dbEM[NjEEaB2__HM_eRo^IYSY90^_1EGEN1DNbgNMCZDYhi
@;gG`:KB@PbiEb`FSK\<\HEmaEaB2__HMQ]YVO0bHHLGkOSGUjBR@l;6E@Xfjk=p
kUB0X0U0Vk?`CKcGEg3nLFF@E=g_k;Y;le>Gnd\k0C1G7XoPE28gS80A5mgYdHIN
k4;;=8Gh`6>cmKcCEg3ni\<;S=g9k;Y;le>Gnd\k0`0G4_kGa@>3Gb3HJ=F\:8g9
f?;f=8GhVk>9mJKo^^n3_>F:EiJ[5UGf6=cJM4dnX2Ng7FkTa@>3Gb3HJ=F\>W3G
TG8<dGUG5PV7AT@SoBpNEkcW38fhULK0@;IKQ2@nM4c@@o3E2=0^bW\L16:g6e<@
:F_[XnCDTToaj\j1lJdpmdlf8ZQWMnilUSdDoDNiMc:4<fO7KD]cXQ^LgcR4@jmo
mGXIDOa;V_XLKlEjIEdSmcBDfFQ;M1PT@JdmoDNiMi<?W?T<KD]cXQ^LgcR4@jio
gC]jnJ0FgPG4\^6HeUT:72IX]ZVmK@i;UUNI]H8Qh7:5<mB\_J2M75DM<4aGMMYe
lGWYEJ0fgPG4\^6HeUT:7F6;YO`4:6iH;e[AggqSn[D:kdYNmH@kgWV=8HB6MTW_
FlLlV8Mo6OmYPJ?dN2jE8E>L100DbNe;@KkMm08S6Dl5[dcNm[@YKWdE8Hn6MlWB
S;::38ko6OmYPJ?dN2jmkcARoLiHc36TSG;E6UDBmQ?5[dcE1Z<kg30RJbBNL`k;
FlMXnXa3>2c9CShnlGVVIEk;gLoHc36TSG;E6UDB]Sief]DN6@b]j0<UEp73n`K`
>G\oPV4J[O9?X9H@JG>_<k?[4<0mZUnY72`oINMf>WYBkB<ZEX0C?N8_:A?mb?;G
>:\oPV4oc:?me0S@J=>AR@;`PF]4ZAnY72`oINMfVW_OFlYjNcF=LFMR>=SmbS;G
>:\oIV>1[C9=]<Am6U]DM6?[4<832bceR[=^PJAlmMHZFeYjNcF=LFMR>=S<0FRh
RaofTme<XSdBqfOJcTn`oKo5KJTcR>ALd4C^m79@DDL8K9S7E:OU?lKSK[RJSfAJ
O<YXHha2cTL?WPORHB0`6Ko5KJTcR`@<WB0K^=F@]DIXLG?7J:OU?lKSK[RJSfZ=
XBUD=VohjLL?WPORHB0`6Ko5KJT:i>7L74CL@@?:T\4[e9SkJPoRnF:?S\OLM85=
FBUD=VohjLL?WP<;Jo@Oh:7d09HQZdKq0\ilVIK@TcbHcmLIUj;T0[7B0QbC`Pdb
hQb`KUnh?0QlFU3c<_FNUkmf[^[WcYfnQU1gMjK@TcbHcmLIUj;T=i@f<45o\5Q?
WaZk0Qnl?0QlFU3c<V0T:89C\[[lcYfnQU1gMjK@TcbHcmLIU=EAgT7H0QbC`Pdb
hQb`KlR<SSD2GA>mjf07:89C\[[lcYfnQ_k4Fai;iaBOPRY[a]pHV75c1dh4`D;2
:76RZijQdY?\D383o`\U=7lf3BXi2?kbgCWaCnRQ>WVYDI?3hK064AW51dk4`D;2
:76RZijQdY?_6VCdlnLGd2cF0`Ni2?kbgCWa^l:6VZ3YDI?3hK064AW51dk4`D;2
:76RZijZc?Y]YjQVo`IU=7lfNXLj_PcQJnl1Pl@6VZ3YDI?3hK06;gERKSK5oLSk
?ABC2qG9WS:Xa_Io[BiQn0aX`46ki;>:<G0^O4`KTH9kZRX8NjRa0NiDkX[533>Q
40DT8he279M<a:Io[BiQn0aX`46ki;>:<G0^O4U@WS>Cf;87NeRa0Nm=^A7Q3=>Q
40DT8he279M<a:Io[BiQn0aX`468YChAOhFeaPaYT\9kZRX`<WffjAei^]7Q3=>Q
40DT8heMo`2e_I?E_8^BM0ijp;YS8>hIFi4FBI>l6=eW_;P7fo44_9jET4_\8LDa
fP`P\068XNETNajTeFNhMlB]]SPmb]RIbi4FBI>l6=eW_;P7fo44_9jET4_\8\V_
M:ePO06KHZ[3MajTEFNhMlB]]SPmb]RIbi4FBI>l6=eW_;PZ]F?LVo6Mg98bZH:>
=aLedYFQhZ[3MajTEFNhMlB]]S=U1VFUhK[n\Ma^Sj1pVS;2SQI<nG^;G:6NPF[6
Pc[_?D[E\Col;7qlI_8<<@VDR<6JU_1O6T]SPQKi>O@`[aORcn@`=CaEdPlCX72D
H6D[\B65];:5<1SS>l;EK@VDR<6JU_1O6T]SPQKi>O@`[aORcn@`=CaEdPlA=Oed
KK`[\B65];:5<1SS>l;EK@VDR<6JU_1O6T]SPQKUaH4`@G22GF`G8\SEdPKC=Oed
KK`[\B65];:5<1SSm[WU:cF@g6iCkUd\cq^\Ma99:5K0f;YB5HYUP0QLVV1Iih=B
HAD>Og<EH43WTAFmDdjgmg[XYFHjl4CCn<8=Sk6D:cK0f;YB5HYUP0QLVV1Iih=B
HAD>Og<EH43WTAJbamRgm1[XYFHjl4CCn<8=Sk6D:cK0f;YB5HYUP0QLVV1MZXO5
[KWEKB21S;hWTSJbamRgm1[XYFHjl4CCn<8O4k96off4iI8fciQ^pD8n<\[N@^f3
]hW_@OYdN14C`25A443ISB:3kZkT_SEg06N:Q`4C9KEia0>;0h_:?WQK;A_N7^f3
]hW_@OYdN14C`25A443ISB:3kZkT_SEkj]8X1^4C7KEia0>;0h_:?WQK;A_N7^f3
]hW_@OYdN14C`25DH5bJ_n:3hZkT_SEkj]8X1^4C7KEia0>;0h_:?WIaBE5eRg3>
O>MXTLHq`DX]>87_il[L?4NoEDWA@\l>[K;_kGcb_X46]>?;707kJ32;_<ohI_BI
N<Om?iaFk<JX;b7Hil[L?4NoEDWA@\l>[K;_kGcb_X46]>?;73J9lTEX_<ohI_BI
N<Om?iaFk<JX;b7Hil[L?4NoEDWA@\l>[K;_QX`[b]43]>?;73J9lTEX_<ohI_BI
N<Om?iaFki3TMmdYG1E4LV]LO1p3ZnF[P@YcMWNde=^^^Q7[^m[WPRUeNpbf@YDo
S6GfSdS4daYYXHIA\o`05PFSGgFNB?olb5RaYG<SSA]i5khF5lAgn7W5U7fXTgPR
S6GfSdS4daYYXHIA\o`05PFSGgFNB?olb5KRg]T\S>]i5khF5lAgn7W5U7fXTgPR
S6GfSdS4daYYXHIA\o`05PFFoTZ>j2olb5KRg]T\S>]i5khF5lAgn7W5U7fGg1QY
VBV2IDbPD?O4pX`^6?TdY^YJoXX4B>4FEb_[FOBI:=_\>Lnm=P^gn<RiPhQAeMOA
L\fV0j50PF[kaSMXF?o^D0f]i\l?]^EFHb_[FOBI:=_\>Lnm=P^gnKEdTd7A5MOA
L\fV0j50PF[kaSMXF?odi^YJoXX4B>4FEb_[FOBI:=Q9X8HW^Q^g8KEdTd7A5MOA
L\fV0j50PF[kaSO5\0R2X2aW_7nlF;opWeD;lFPKo;j803AdjO7C;[WgDFIeKKOd
^Sag2IFe[;392=_c2EB_=RLG43`X_]eof8nQJc64<[bmRNnOjOeai[WlDFIeKKOd
^Sag2IO\[mail=__2EB_=RLG43`X_]eof8nQjKPeo;j803AdjO7C;[WgDFIeK0aX
AECa^IO<[mail=__2EB_=RLG43`X_]eofeWN;Tm@K`Se<@4>L4pSZJ2UJ6L18>M_
MABWGIX?YPmPV>I2MA`hNmM^Kcf_8C0^@UQ:DooUfjjX8E^d0eYaEQ>=YKcJnU4\
LfN6WKogIPVPV>I2MA`hNmM^[JKBP[D^@UQ:DooUfjjX8c6\`DT6VEI>36i18>M_
MABWGIX?YPmPV>I2M0dFMc:?[JGBP[D^@UQ:DooUfjjX8E^d0eYa3XN3f[iEGMCF
9Z4aoq@Ee=4Ij=1IO83fAQW68S_nX[W^aFeM`k_V@@^CdU61h7jgc?2]ohjOnYM8
ECMf;H@XhEPI1_;POP3T0V\ZF9MeX[W^aFeM`k_V@@^[ElcT58jgc?2]ohjOe?MB
VffOK^@XfLiSjU1IO83fAQW68S_nX[W^aFeM`kQVBP;DEUcT58jgc?2]ohjOnYM8
ECMdKiUbCOZ^0BLMlk6OC`4oqIIY5JP;_jQHSjAAlMec9j;>@MO4FhmPZ<=`JRHS
VpPa`kQ4F5MLMMG_TKBZ9<4fKfLkFHiXAldl_SLE[[2lYP^G61;BTR3iP8MSCN3H
`aPeHVBN:>f>C5IO1JOLMh4fKMLkFHiXAldl_SLIh@4V9d^G61;BTR3iD8=4M^6E
`?PeHVBN:>GLMMG_TKBZ9<4fKfLkFHiXAl1cAYS[h44V9d^G61;BTR3iP8MSCNIk
=2\RPTUa[goTRoXi@jDSpSPnEh@^[Vb\A3RW=B7;nLZd`N^@jWAnYK_;0QRjSg1k
N?Td432\E7?c<XJ5JQGmGSk2FZJ7h]RToE<A`amAXYZd`N^@jWAnYK_;0Q1hXl9I
<?Td432\E7gAQ83o06GmnSk2FZJ7h]_\]3RW=B7;nLZd`N^@jWAnY4B^lgfh=l9I
<?Td432\E7?c<XJ5JaeEI6P4Faf<R^1D_cW@bh^qAaL`AibXj^>=l:IJ1hBMZU?_
ZQYGgXdQkT6>>>l0^ASUUSJR@Pm`dnS=?39Ma>4OA^gP4@MIQ@DQddC2G;BnZU?_
ZQYGgXdQkT6>>Yfmf48YUSJR@Pm`dbYU:Ra1<>4FA^gP4@MIQ@bQ0:In1hBMZU?_
ZQYGgXdQW7=V\ifef48YUSJR@Pm`dnS=?39MUFVjVbdL]Fo`FUD1Fjhc6JqQ[E<n
SB49]d8jDn1jE_C0OjR[25\^A2BOL04KF84oWX_[k\8ZleDgZ_QMO;7gIe\Q:AR\
LiA2[>=^=@Ehd_=0OjR[25\^A2BOL04K]O\]oFC[k\8ZleDgF6WNf8^1OeDQ:AR\
LiA2[>=`VnjjE_C0OjR[25\^A2BokJ8ElOS]oFC[k\8ZleDgZ_QMO;7SVigSK_69
[BOaD9LcFmBnCp6g8ka5\ghLe6_IWXV0En>:^nP3jm0c72QSCdieCbdLEXL3a\7j
9U7m>Zk0b8bai?To=]Jmd\24]a6<b^V0En>:^nP3jm0c72QSCdi<obc3U<L3a\7j
9U7mXoC4JQBYa16o=]Jmd\24]a;\W\V0En>:^nP3jm0c72;EiM3<oLc3U<L3a\7j
9U7m>Zk0b8baIl_[oeX9IKYfj`\6fGdoqPZkQRSYQJKh\f>jJOA\fA7``:b1hFc2
Ea=3i5J?Ri[6V67=K<>I5KXk9e9mYe5Q6e<b3K:_>[=khf>jJOA\fA7``:b\LAo0
6>c:33SK]i[AV67=K<>I5KXL9JVE_Oh6<P>l=CMeGV37E:mjNOA\fA7``:b1hFc>
\>c:3IA\f7KAK67=K<>I5KXk9e9mYe5Q6ebhO28^TaH^0j[0XThp7GcnSQB>PDZ_
mAi@l<]]KJ0PZ^_hmK;hj^J;e0DLm\ZYk;f63khb?<l5iET7RFE?fe926NB`PDZ_
mAi@l<]]KJ0PZ<\Wl7QZ;RX:^SLem\ZY3IfI3khb?<l5i6>7Vl`n7fQNc?>A0Z9d
c9i:l<]]KJ0PZ^_hmK@h;RX:U9^]bncOY;fd3khb?<l5iET7RFE?f]D>Gk_bm3N;
jYC^TWq=C0SHKK`jZXbGETk4P@R`=GYFgITD2mhM01iGa81@HH4bAflVo`HUO\k;
cehYV@aJd6gW6K@jZXbGETk4P@R`=GYFgnT[f\I[k1BGa81@HH4i>kKVo`HUO\k;
FfL464K=>1l@PN5nS<;VETW4P@R`=GYFg?Tg<\8[k1BGa81SWHK=[fAVo`HUO\k;
cehYV@aJnYgcQZQU[c4^oRKXbq\93B\b>OKS3<9;IRc;YEMLce7UhJEJ69LK2>gT
XICcRbFLWTJQIj=6R`2U;nHk87JZHH=_>lKS3<9;IRc;YEMLce7UhJ^i6bLK2>gT
XICcRbODNT;VYK=6R`2U;nHJ2P5;:=M@b`lS3=9;IRc;YEMln79VZ^6i69LK2>gT
XICcRbF1N`;VYK=6R`2U;nHk87JeZSI[C]MLi4C6hXP6q1o<Cf;R2GbnC[:;5eZW
1UiALVQIYij:oYiU]>Y]JIi`^1OdaCThg]MQc?;pI^lR9_D8Wj>o7j8K4bZ_E_4o
\jEEPdZBe=bF?8G>T0XbG\XRW6Q:M3H>mTn?Ib_IFKL;l?DMWj>o7j8K4bZ_E_4o
\jeE_85K5=bC?8G>9MeWT6W`hLgV]PHImTn?Ib_IFKL;l?DMWj>o7j8K4bZ_EfaH
b7BJ>dZ5e=bF?8G>T0XbG\lRDLgV]PHImTn?Ib_IFf3c_kULjN7i[FkW>Cq6Jd^k
A>8Ra6ok42`8;Id;cVGhgobm3in5eGUHc:Mf9J<ST;V:=o50XIIG5lRFC:2]CeAT
U=n06n`a42<nHeY;cVGhg;G`79l7?GWlN6GWX54RA;heXmN[WO]a5:56C:d8>g=T
]6K0612k42`8;4JHWZaPUL<n3ig5eGUHc:Mf9J<STfYimh>[W[@7RlM6C:d8:F;1
0[2ZDocK>>DC5pl^b;<8Xj?jkKW\6YlJJK\H?1F5B_PcW73FN7aUnYJG<<d4m3Pe
9\l56ZL5;7WQZSl2g1CGXP?jkKW\6YlJJK\H?1F5B_PcW73FN7aUnYJG<<d4m3Pe
9\l56ZL5;7WQZSl2g1CGXP?jkKW\6YlJJK\H?1F5B_PcW73FN7aUnYJG<<d4m3ce
92l56ZL5;7WQZSl8Bn??K38?6nIZ6_5lqBW`0kRPNM9l]0noX8B2TTg[[^LERLh_
lF[fPMCWF[jhfRT1XJjg27_GV0o_Mi1ABI?oMJ0PNM9l]0noX8B2TTg[[^LRRgmP
DUWD]37IMmiL?=FG<F0KEc;3X]o_ni1ABI?oMJ0PNM9l]0noX8BHTHY349eU=Kh_
lF[fPMCWF[jhf@FGXF0KEc;3X]o_ni1ABIIf2aO^?mnKRDij1ZEqiC>jFX9n94NA
fC;bXhdbd8I3eIRRGC[68MH8Q8H8C1\a2;;6C2Fo@bhH4D]9S6TlU_;e:=9A94NA
fC;bXhdbd8I3eIRRGPGh6JO9?;]JMYjL91kTZnho5S3A4D]9S6TlU_;e:=9A94NA
fC;bXhdbDTQ`Q5TekF[Q8MH8Q8H886oW91kTZnho5S3A4D]9S6TlUOn6DR8E;Kd8
XMK\@SpQjOg]CAQ\fV0j50PF[kaSMXF?odi^YiKOe7dYMGDj?TDYeF<5?\1Lnm=P
^gnKEdTd7A5MOAL\fV0j50PF[kaSMXF?odi^YJoXX4B>4FEb_[FOBI:=_\>Lnm=P
^gnKEdTd7A5MOAL\fV0j50PF[kaSMUV5YjN<8]5\l?]fEFWb_[FOBI:=_\>Lnm=P
^gnKEdTdLM:Yl3cGB;WRf[Cb0pX]m^ibHHWlO;8iKS38IL13Y?bBe9hCU7hoZX4:
W462N8G;YHTnIllAKMY_F`l[gm@0Q8G]HlWlO;8iKS38IL13Y?bBe9hCU7hoZX4:
W46;O8G;YHTnIllAKMY_F`l[gm@0Q8G]HlWlO;8iKS38IL13Y?bBVnmG5_hoZX4:
W46;O8G;YHTnIllAKMY_F`l[gm@N\OBPMTc>^XgH<[V;pMnDHWZ3QF6<YNT@`5jb
jJ?GAJXbFmRZ5\1eq==3W3LBqnIk7kaD$
`endprotected

endmodule
