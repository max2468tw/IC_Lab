//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2018 ICLAB Spring Course
//   Lab05	    : Workstation Logging Simulation
//   Author         : Ning-Kai Yang 
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`ifdef RTL
        `timescale 1ns/10ps
        `include "WLS.v"
        `define CYCLE_TIME 15.0
        `define DELAY 0
`endif
`ifdef GATE
        `timescale 1ns/1ps
        `include "WLS_SYN.v"
        `define CYCLE_TIME 15.0
        `define DELAY 0
`endif

module PATTERN(
        // input signals
        clk,
        rst_n,
        in_valid,
        in_data,
        action,
    // output signals
        out_valid,
        out_data,
        out_action
);

//================================================================
//   INPUT AND OUTPUT DECLARATION
//================================================================
output reg clk;
output reg rst_n;
output reg in_valid;
output reg [1:0] action;
output reg [7:0] in_data;
input out_valid, out_action;
input [7:0] out_data;
`protected
IAYYXSQd5DT^<hPHC47l2ifamiAmo^afTA2FhjK>C7S2<ld[Y6pW_QFT]F1_0QP2
gLDek9abe=UVg6kUNZgP9SfD8K6b8Z`QOgqjA3Q`]1`LFC70f9G;A9epdSVk0cqR
MkkkiO:W59A1UJ666\M2]mGcWd@H9K?ZHSpM^NFL@\AEbJUbUE17U1XkClacQa@q
Yb\n6NbRn;ml`05L7TeVf=mH@=q:FjC_5MRUk`hamj6JiO[_^SE>AZ3gD0J7ZoIX
9ZfdJGlgeVH?k0pO11JOVA^4MRC9E51^?V0E<2kqkPNHJ;2GE3M_ngX4_P>Xp>Jo
LIQF2oPmBW;9ck:h?V6q]`FC>j\5IEH=IPj;lPHfHUF1O:nkLED=00L]E[PSF7pc
ID1J2?U]AlB=eS[Cif72l0IFHXBl\WM;XH1?Qh@=V6dJV]CfWOWTlV^Gi>9]]@7p
oGDeo<gC7M[JD:31V2B?WgU[]M@Yoh3nH=[kpKJEY?Oo\hIFaC`@SR64ojNS;n7a
Djned4D`jo8cjHgd5goQGF\SqU@c[k3T9TNlNlUF9Ci06Y;^\mdRU]S8dXFD=\oT
NZ5C@9JMi9mcpLC:8aHi1<b=i4l9CS_D=ATSUWYU3qRBIS?Tbg<kL:2I8H29K?9=
=:ochME>_4CIlg6M@>K55F77NG_=VVq?2o1\A6aDg22P@kVh@>=<\^C>5ReQC7b6
6pTh3cUKAcIFF\D>[RF8T7O2^73jclal1QK`a`mQGoWDIO]Pp:eE`7ec`iS@Ya\f
<;3eg>DqR0MRUWY9qDHT7S1[<`GdM_1SFVc=qUT]WCQWe05<;mR8YV8TPn@Blj?c
ep7eJR0b8BR3abkjJN\`5I9=V<4YfCO9l\qQV>`cOh]F;OLlnD7DI\6@a7j5DHPh
Hip6d[Kh;Sm[=5@S<L<@lI>j2gB^hLkI4p^gSeV]YJ>9A;WnK>YLB1K0dpI1T<7O
?TUIW=:]SUHiFbQTMn>o3HL59fZnp=?4Yi[N82KSf4FL\Yc^XPa3gfPgEE0RqK8D
2B=8SQS7U;@]6T>FSM0]\ADMjK\V<^\gTEjQ8<BHlS3UkXlm`YY?oRF8S;j?<UZ9
fZ^Y\_mjXP`1^H:]o;_lQ69^:8VBL>CTmHPE3beffHO[45>f2J[cpk3kWb0Om13H
^:hcT_R3NlCf0[V4VU2^UZK[@GaIp7lAALHE\K6m3RAYMV=ZZKM<c5llR`>BC^n3
E61kVSo\M56q[:Od0Na6O[:MhWF@0EDE7RML9RbIC53bq^H\^A8F7lK>f9UCMW;6
iIcEk]_87<?HAEj[76M21QbWhNoNVYOHi1<`cJ4i5\WTOif6db=kWYdP:`4c3SF1
K<f]7p2^c?jBAkML93WNMl2<UQ^hpaB0CCo\KX7d1G?T5Y`PpaOR];nh92[We132
p8@Ha?B8DN3_Rh2T32EikB]G]IbPpY8F5iUWI;IgcA96Ql5m`pm>;D<ahpN<jKQ^
XV:^3Za:Rm6`\Z_?8O]2p9mQokAYJIJ^H4SXIdNnJThUY<6j=bMe>G\PeDLK:1O_
`3Xa4bN[U``VNUAc7<M>pcg`^L8pDUKJaM@<4V5UB\V\GieIY1Jgd>c<`kL:TPOp
A>@B=?J_0:NVRj@2ae3Khf846j[E;18P<Iqf79?MlZfjgY2FicV7bq[Q9hTl\^=A
oBR6jEoJi429h]@^`7f8VhHI=]43:G<LPC7`B^a[f6_aO@V<NA@7D:oWfYIOQZnG
K_<[M@oLLm0S5UF=XNPnQeHQLg:i\qQJiETW8E3iCUBIaIU1RiRY^8Lgi1M47G=]
=4R;67b0]Qn[:QlSZ4cWK8I4dh_8I7_g6b=W8E3iCUBIaIU1RiRAS?NY9DOoK?[I
ZdTFiq8BXU4=;3hJ^BVj4N=I=cdL<1Wm_E4kZh27LRIGgSZF51@B\CoQbmg^HDlI
0P?nRk8Uc>T9;4hJ^BVj4N=I=c9VKID3cl6HA5cQLPoLeqa6?SX=P@l:mo]`2Bn3
9J^K[@J\4]ol4`N?WQVJ6`WnQDU_O6G07SfcZ_K>8>SOE^U`EBMNa]B?K77L20DX
EP^kYQ`]4>Mc_jlA91N=6l>F:32d6pTLCPg3IdQTmjjeHWJUUb<gIPS`L:fI\;lc
FdKNOa?]PHS6>Sc?KD@Y_]IGbNhE9YpfL7N44mCZ9LH2=]bGBiUVS6CnU:9mc;7>
MbUhlB31^B3hK]imlAc\WC1AoPNb8WmnVBQN4mUZ9LH2=]bGBiUV]QJb2Jo5@5f>
Sd5f\7q=kNiHbKad52Y`QM4qJo_W?JMqBN^MhlZJl1SYO_b2enA8=gL[0cG4d_ce
pKk4QYgjJQaiA:4R\UR9]@OkYk>pGI1]XK]<pX]G[WYkPP:mZLVa?>DLTGli2=Qp
JXb4A_]oNf=GSBan3??6qOCgMigD7Oi:;V1Y9Cdl@W7CF6GOqTJlZPYjNWJa0J1_
CO\HJ\fU6KM=g_`l]pf;f2eSZMX3ck?`j;^K^a;b^fcUjkJO^D]SMO3:C]Xd3?5D
Hd7bmB;gXlPQeSqj]2=m2jd2<8?cn4:_0ac`W^Z^K[MR<XD=;\pWX0KT^R>o]ATD
n_6Bb7TL^4f8Z`M1_6lFB>qmRm5=]k=AQoF8:LQ27=O6lkmPZ:Xn[O12Z8lYid=R
UPLh=pKJXFIDfR>c\WkA\mUR9S73YJ5NPXNTA>X^Tiic4MIaQUMn9A3Kn_gW];U;
S>QXpDdacgcf2[DI_^8La<U@WAL0ckRDqIR6@Ta=T_j<U4>``3koN9@hQdY54]XZ
Yj85;C[:i`f8qmjMUHHDOo`G`YhOiP53pg1Hg3oQKJFB=BZO2\Pq:F1d;o88;^3o
=GARAZJ?\W0foKPW9nq[W1?PFlq4YmVB9b1::pKIBSQIF1?]ndcUm`WVYq^m\8K;
GV5^DKK[\GPho3ffB<Z60SnSq^D\WecGpa_;Y__=XB4145F;U0c]D>F]b3L<[mU:
aRLCq9]?1S2^daX6M;LUh[oMVSibBHjZkT^c?pJWaZPhQHCheV_I9lbFbRF@h@TS
0eW07qdiC;`XW;pJ`cBQ1jW;=I1JZR9a>SHn0bqYF0e8WP:Mn8YI]<W44>@qWIMI
[:[JmeZT=NM5RodS_GZ6YgK3G>K1;:Iq8>L>]LiL1;CPgX7EVf6WI[Leoj\?`1ao
CbY@?\>=KkGkXPADgnf]f=6Ock0O^bpM`^TKc<j;_W2JQZnOA305Q:d`D90WOTPk
enb?UUod8dmSECJL`8Nec;S>cNQZYEd]a`oCg>U`:<<n]HUeli5gYKQ1ORO6kdSS
<IkLnL^@[T3]n6X@UQIj?=Fdn0MU?Vao=1;Q23f?=NLOc?T9J8oFnpF0j]hZ_C3m
WaT>e?TJ03ThI3?`<@cOPH`k<pb0Glhc^VWKF^=35qjd6Nk6_pU`onTKAqUlGEIY
;YL?Ok@]4c]R3eo3OgVHUL=\J4`e>p]bAEgfjT0i?Nh6ZW0kc2:]K>VHNB[jHAR^
G0:kq>Q2kZY=7d2ZH@k>>6lCc4\84GR6e9Gam0nQk9_9io4>iA\SI:KZq2B^o0_C
^I=oQjjHjg234fY?mA`U_SOnZ^UYe92ddfkBDo4Tngl4ZWoAUUb7oo7PiGjUNJKK
3L6NVo77?1hYd79VBCcRK8=RlFE]kY;25<DYU;>ZEcIl3QF1T3CAZU3hICfcCBhJ
IfNIKijKH\7Zg7_jPqR]4=6f[G@_9Lo\ci=5_<OXA=kg09A3jI^Y]6o=3C;MF5jj
]0k0]MpSS3HHPHW17U=1BmCMcePWhiiBPZEe72mNZbpmBlQ1AIpcT_^co1q5;9Zf
HF8hd8C93:X;Om@101VHB9`HVjlkK6pK3@;<SSk7^bbhHnCda]k9XMP?6ib[D=?8
9@4>E5Qp=:=nRac7DIj<oVgYB[?fo4T8nGRdQ8Jf8h[pKgBoTIeK3h5SHe`B`D5I
;4UbSh3SHMYLC;U4?LT@^\BHPT_p5>7[l1SC18Kf3aKAdOdMNdRBe?Bj7O8YOAHF
eR==\6hmM[d[SF<Uo`2ei<a92?F;hnYp8JB549CS1aQmk0WU^gNKo[>R?3]FDUPh
Aol\4mV^Z_Y>Q1nb:1@>f]>`0BQ805^p[:8@C>\XlXHRCf7Y4jICnGG^g5GdR1pl
7gCEXKp5<XkeN5KTG5Cg>8M:ODS;Bomkf^SAjj6k3a0F:kSRC_]?2E]cP2pfWf5f
FapndITneK?T6K^7@kck4SFiW6<g72jnIQQJbR1E61peb`omL:Lb>Q5R?8@?QW9U
VEK:;^>nkVa?:O<R9QI;ZDdUn[eAo<0b@]mMYJ1BlpUEDEi_I27S;bc?CSPIm77_
WhIijocf?cbS9UQS<kZ\Gb8__G7Zg;]i:om_q>Q5d47eBj=fN`>j^<?OH>FA]4@Y
ZH<qB@E9T:Rp`2^<DD=pRdfYSf<fh1CJ0A^aQ@?ge6J@:b3W9_?Z^3_0lRJp61j7
Wm2031<]hY?]N8CDm=:KRF9W6kbiQSBAQP9NiUb<XJL?oO5eq7I^ML70;E<kAdAP
1B5\MmACS\fbOC^Lbe[\8\@cB]1m0aE]SlD2iG_X_SRPVA6W>\hNqIME?bVMSe2a
aRWF:n2BaP7Q2;8IOm\L=3T5_`a2Km<Id8eWAhEQDYG2i8cjQ;kUpQK7DI\9lobN
YCBM?SEY>387=aM7\LRqE3Id\gIqFd_6dEAd688C2@Tgqd^CldeQqJ287LbLL?id
O>M^JHBLZ`ZbYfLoXh=0N2lMFZHjpS]gJO9lpRCFL;95PTmpnVeCL?ba6`dX\CA7
SZJN4Kc0C6kj^A7CIIiSY]\naL<nLdqBVRlK9Z?FlGNP^1fd\E7;=TGABZSmVZGp
63RWX3kIib8Cm6Q?9K3A7?gPA3`MTh0Ii\hp2DIUQJ>DiEQm9mCC_1i8`AXP=E[T
4S=J[;<pH48oDk0pIOL\L9oSp]0B`foo10C`oa[>2fVGe8V=T<\8K_l[p@R=]3hW
B]CIXYS?NBlZEV6qj^7l:WJ4gUZ4TBbW`F]]:4;M8[^_a8FiPCq\=X:TX07?egXN
OC=A_k:j[adMO0NZ7p`ToC5L41I5jnUnhmnlH_9:92SMT9qX^J?ioNG0PK<9l\Pn
oYRB2Jmg[_5LRC;mP`7WDgh7IiSiL06FGXR0KhW;3n]o_C11A@3?oNG0PK<9l\Pn
oYRB2JmgaJP6jCC?fiZJloS3@Jq?g@31^oN?A^:?ZNkPLH_cSqR=^o;;CMn[4JJ9
h4Gh196[_hCGZm;6?I]cQhhkX8QDG^_EFfK0^FlnFEChYWX>TlRc^OJbC0n[4JJ9
h4Gh196[_hbRFF7?6bSBC[c0X8LKfpii2@5Odc8gWY3XhXV6l\cB]R[YOX79F_F7
Pm2dcG:V8oP`iYHd?8iEGj[X]ETcFX1kcm?7dT?Xl63XhXV6l\]>1^?dD;1=N;40
]E8[T7FLZpJmS=4NUZD2I0gV_ATKC^35VPIl3]`2BXBf3OCD3mX9F\LS56?CJ_g0
b?:8e2H][cjCc50NUZD2I0gV_ATKC^35VPI_oJ5EElZNV?=:_Ig@1q@WbY0O7;k>
LlDUKFW]g`a>lh>LkOJ0b>VNT1Ok_mei?=3^d0]LQmX?p6fRTcRUT7\iK4J<R`8X
8<RN\QB<ql_mJ[nHjfLF7hm>cp:IiJG6<p>0H5ToaLC2hPIDEW7=;q0BBJ8MD?2`
6i6Va^:S=b;f3I_7@nEdfNbKf5pRgX<?><poXX`lb25F4[l21P]Yck`1>TkFT8jI
Z29fg@IGMm^Oe6]CDU\[UYV]6ldHnpl4TIJo2nq68J?]0eBQUa0eZHdnPR09JhDq
odm;_AFlIW8fao3n2Vq[]<__7Y\E\=8XT[kjYKT_[7@VnbMnh7OUnSg00j8>d[=B
WLDNGVo]DWAcAp>;kMU8aeg1Lc0II[bFHkJG2q=NK1`6405TR@TJSN_Cfe>O\e@g
qbG=5:_Q7kVghec[hCaRiRD[3R<:l2?ITiTUMYDqbh@iB31]V68\:K[X9\lq[\Y4
F\o;^VQnZV4ck4[7e3FSL=iIbRZMG]]6pNPJG[Q4FZhR0W?9XUC5>Ch8e55X;U;S
EVXRY>RnaY1P_86;P_N9gLZ;hRj\=4Dn=hg4f??49ZhR0W?9XUC5>Ch8e55X;U;S
EVXRY>RnaY1P_86;P_N9gLZ;hRj\=4Dn=hg4f??49ZhR0W?9XUC5>Ch8e55X;U;S
EVXRY>RnaY1P_86;P_N9gLZ;hRj\=4Dn=hNHHjPH@72>_6O:P8QBNq0@F]7>M76R
`aEjEZX1?]3o6@H98Z2H:j<aL=]YHEBNET347P_E`4A>1LH;E2gC_M021;Y>M76R
`aEjEZX1?]3L62Teo>Lf=4jWa<SYHCBNET347P_E`4A>1LH;E2gC_M021;Y>M76R
`aEjEZX1?]3o6@H98Z2H:j<aL=]YHEBNET347P_E`4A>1LH;E2gC_M@S1n@:K]_b
KhiPEWZ8PpWc3jcn6Yj_O@nLcY0n?@ADQa\CYlLFK5^9AhUolRmTGWE@`GjG>E:m
_<3;ESEJBIW>aT4\NEd_a3nLnYhdKc`@QRBeYZDFUhU9JcWFm<m5QFEAZV>7jT28
SF3;ESEJBIW>aT4\NEd_a3nLcY0n?@ADQa\CYlLFK5^9AhUolRmTGWE@`GjG>E:m
_<3;ESEJBIW>aT4\KA>_3C8oW]<RU@PDCifmq7LL6J>[GIW=P?hdifJ\F4MO\glV
]gFl^LVin;B\RT:5[Hh<FU@F]@n<Si>]LdX;Q@BLKP>[:IW=P?hdifJ\F4MO\glV
]gFl^LVin;B\RT:5[Hh<FU@F]@n<Si>]LdX;Q@BLKP>[:IW=P?hdifJ\F4MO\glV
]gFl^LVin;B\RT:5[Hh<FU@F]@n<Si>]LdX;QU4D_515]o5cKiPH07kmpUdUF[E1
VUMEU?S`XO^W6mgULJ47^?HLaq54gP9<3JM7f\^51O7R3cnaiVF1a^qF5RmQ7eKF
PVnW?QQp0F`J?:7qRV1H?T>`ohQ3J<gknTD97=mplB9oeAnF;^e@Df20jH@]B>P\
HQRqcd@ES;Gm[@`b=lda1V=lHC[gTaXBWo17Md9>;IAN8S?F_mF@dgeZN8GEK>HU
Zj\of_odm]G5[@`b=lda1V=lHC[gTaXBWo17Md9>;IAN8S?F_mF@dgeZN8GEK>HU
Zj\of_odm]G5[@`b=lda1V=lHC[gTaXBWo17Md9>;IAN8S?F_mF@dgeZN8GEK>HU
Zj\ofA]a9JBbjQh4QiN:iNT:p9[Q35k9`KC^`YVY:5NT3`AKOb`Nhe^PCC`bdDkS
ij]n[?=LWe0k33bCI];4OGV_d9HO3\k96KC^`YVY:5NT3`FKCmcBOYDGAoLH3?kS
mj]n[?=LWe0k33bCI];4OGV_d9HO3\k96KC^`YVY:5NT3`AKOb`Nhe^PCC`bdDkS
ij]n[?=LWe0k33bCI];4OGV_dYjO4<XoOk3F6ahM?V;4pbM9fZ]8GlahXbXAYN71
k\[L]VClI\XDSiS<fioZ`BTQ8]DV8dMG2G1@<GHBD5JJLbJJBL62dC?LIbX906cj
:oOLF\flI>ZD\>S\`g\:_B6cn]6<RFZ[;K_5jGHBD5JJLbJJBL62dC?LIbXAYN71
k\[L]VClI\XDSiS<fioZ`BTQ8]DV8dMG2G1@<GHBD5JJLbJJBL6Jbd?<B_b59^Sf
cW<dn8VpeEGOWi?oeCn>2O3MBN;VGd>MZYBc9a9JCQ<6a1a;lG2Pm`0XD@][e`a\
BH5T<ed=lZfGVi?oeCn>2O3MBN;VGd>MZYBc9a9JCQ<6a1a;lG2Pm`0XD@][e`a\
BH5T<ed=lZfGVi?oeCn>2O3MBN;VGd>MZYBc9a9JCQ<6a1a;lG2Pm`0XD@][e`a\
BH5T<ed=1_m;9lg9iALXVN?oR=cpB:0?5PQI_[MR3RXQ;SH>`9UOB\M:D[TY?od?
L[mie[dn;YPAf9VH`\=jD]\pecgAC]W4HS8kEPjDlg6E[iR[TZ\lp<0nnmKF5`oS
UhTA>p[kUK=0agpc;S1jBOdh<=@KniF^BM9`8[j?Xfggm\Jdi3mB9BPKILlpBR0_
makE]39IHCVEl0oQhEJ05FG<3iO]CMIGj]2`Z7cG2N1G@?pQToa4KBZY><FLO039
oSC;CnWL1R5NMKO;K<79NK<gmUc]@HK^oJmn<I_BF?08Ge_`]Nd8aB;Y><FLO039
oSC;CnWL1BTSe]kQBfdXcnNQl0Eq<S4mL38<>G;=A9hCMf37\mfJ\d;mKg4d[]m4
m3KPbVRDDQ:^B;VgPE9K6LPV<kF0<`\^Z[84>G;=A9hCMf37\mfJ\ZP<clHE3J1X
9kSVj1<Yq1nHS>CU4inMbDnJi<L`>G]gQ?Xfog5VPDfD:@:H3:Hi^@\e@b4_3gK^
T9faTc@<I4D4=b;jeinMbDnJi<L`>GIgaP3an>Xc04E_GmmoTWO;JqS[O=O9IM8b
ighD@a`_kN2gEWD]b?h:DO0JH:A?ZQf`979A2XNA@\RIQ8T2a\AZVlS78Fi8=3Gb
5dhSOZ6SfBjgEG2EK42DDahgW5Mo`=mhEL]W^f<h=I7R<9T2a\AZVlS78F?W7>GH
:B0k@2EP=Gi\]oCl:3p0bJFG\Joa_XkQ3GFT`F>IB9hc^E3<=AA>mf4gB@8`cnA1
g=AD<6\^beUIBC23A4;iYX``eJ`a_XkQ3GFT`F>IB9hc^L6LDJQBl[8o9?D_1@cp
9G3g_Z29>8ac33LKFG[\KZMG]?gmb7qNmjPQlY:==dDYQG7W6cmCgle8CJE67p^0
hJ51D;^?=H;N8LjIp3e<4W[Up=b@aagapSKY1Wam]1OBcJAUE^R`nAkEp=CT:7WW
9l3Qihj3I9ZcjoFY?TZDNScS2f^cObCfRngaKj=m_GKD7XD[L[8ep?KTISmUQHbi
hW`e4:;YcV1@IofOLAAghBb\J;=YG9ACf08KCB?jKKhG6EU^Ail\ZiS\kf5PD<?m
>JZI7EG9hFh@N3?4cIBn44=;54OoTfCq=8BCIDTL`G2Xkc[@S[99m;k>Q=DGA]Mc
cL;WlW^Wg^@?T`2V]`pONb`bb?^m0dTOna55RN6i40cA`TZGbT`d`ETe:46]AcR_
KUQMR47lQodKUn3>Ndh<RK5`[?_m0dTOna55RN6i40cA`PZ?E[o]=eDJ\5fHQ?jq
l\Vl:Xm<h[DenUnBp^JMh13CRPHZO;[5Q<_n]cWPaoW9MHblV2mFN>`MG[J^i=_c
KN9=X6D<^cNZZOCmj^h5J4l8VPHZO;[5Q<_n]cWPao@S\DH0=<5I]]R`kDkU]p5;
2fkC:G0]E^c<dk>nB9N8\ThmCQ9?RD@n;K8T23`7M\fV:o1X1XVoFIC2;o]dA?DM
YZ[fPA0]E^c<dk>nB9NQ\5VKkiNGBJiH[9ZC5A5<THp28QWUAfFeB]=lADWnB>hK
c2j=cNmDd?>V[UR>3W:l;AcSleSAURT7\i0A`8oB;7L2:W0i=_8lDiUQXO]@CW5V
G;RKdbo4C[khXZ12NHcK\FG7fWD4RCUjkXSg`8oB;7L2:W0iNk_oDJo4L_T_1RjX
@1U4WUCPcqU09WD^JLjc:UWA<ZA4]@?5ggdH`\g>A^QgiQVGZS=F@\a]AO`hUb>?
f9Z=Be3Xnko:X6H^J2jc:UWA<ZA4]@?5ggdHL\41;UdPA6]89NKZ:4qJGaQYGROn
EOmoEXh]hQjEQU6W:\TPcq\ccL6TRhFQDk\8dA1<FeMN[_8;UB?KDRHiXaOdYlXH
m[1[PPm[;qYg?c\7D8;NR9X4Ykq3?M@WhSqK_QYlaY5[;QK\MKJ4I0GJO5odUYiH
6Xd<TdC:7mXedp\aZC;L?AO[:LKJa9k=8>II_4h1Q]1m1j]AV6nTZYToT=e?S1>m
qP[jD6GMQiH<77oFGh?BR\Vhf@h1_W71o`HKPddD6QJMh`cLFBA^<Yd9e8Z^YG<^
0@egcDJMCiH<77oFGh?BR\Vhf@hkL:fQhC]o0M>ie>1b@pK>Ea_56PjQ:DJ\L]G2
[h`^=aiShg72]N=E:9IoDNM7mc8VkA[_j>2gS=ioU_0@McKNfFm1OkjQ:DJ\L]G2
[h`^=aiKFCLIKFl[cB`SY?cf18p[<P<GY42F_4aYB?h9jco2Sc]KE>A=8i;27iW_
]?kSSl4nQgh]?lOW6PZ]IMqZE@F3m:fKTH3^Pk^Q8iAEOUR0C0Zn?7BO=keb`25V
;mdRaaKceGEY18>:8E28Vi9HCmANKD7KTH3^Pk^Q8iAEOUR`8Ub^ALgFPk\bO9WF
cEbqOgRdclH]\AVIFIdmdaf=O_MCTd5\TFjGVOYZD3\ZoX@GU_XeAcd7`lLFkBZ<
5idfOTG2VJm^TVkcmP1BfcZTBA<XXZG<M^3=l6JAcABN^46RSNj>diM?:JYcSBZS
5idfOTG2Vfi^>V4NmgaYKi\d\Lg7KXVolYqLD4QMJg\BUk\eEK7d7@]Ta4g0OO3`
bA8Q@;Oi866JiI4Pj`G=hk[SM`@[PL`QeAIAb\6VaggBUk\eEK7d7@]Ta4g0OGdm
]DV]LU[noCiXaVMq54F7582>BB^UC62IeUlhh`M4AZDW9<q^5<i3AcTYPcgNA[kq
7`T\K?k<PRSXQ]D36`f3NcfH\AMcm5D16i\b^WCJd@2XAD;f2LphT912e=p72_0G
EP;nICU```VMN8KEm2>1lg\lNog34c2<>[KXaqX1CBG@f;?oCJ]UW9=FFN[<9l9:
LnD9XI64jCWKKJnlQabD6O[IpenVidPeZ<PCdVCgD^:\`oU[D34nFIcCZWX;UmA2
13mh\=Mh]Z]\?cf_f@^Um4mCO4PE0q6oUIPQ:9G2RW:j_G49\lhP]HMZdg>bMB1I
AN0gUiWm;N@AhMMcK@MTkMV_?\C3S5mUn0I6:6G2RW:j_G49\lhP]HMZm49]A2lg
4hgh_X1DRZqC`cUSMXi3`587DLoTf>nHfai_ZOiB0UT527U:n@>ibjFnT0F@i6YB
a=?gU9BM5R@CAK4b31c3`587DLoTf>nHfai_7A;KeWN:MAH74bg>5WQpW:^]BMZ^
2O4:8k42bcL\1WY8a:bh:Gk\8\:gbX[0GW57KGjKWPMZdRO^=HZL4g\6MVfGhZXj
2O4:8k42bcL\1WY8DcTZ^8QI3Y:2bV6HW2hap^d`WgVRECEWT`U0g17gn<fZm72E
]c_V8iZZ707PcX1CLReQO4OKGgVG>UB?GhSMZ^Sn7jgaGIh5g3DZg[6>\9o?_Fh?
4Rd\bc0BmXR<HFMMZAmVEK9ae?W7>GB?GhSMZ^Sn7jI_Z8hYI:YRoY7aiP7NaER4
f8@q0Nni>?6mb90NYei0VPGiAC2DnVF2J1k6T2I438JY41\\h7jZjYDaq_<EB`X>
OlHZbZQ3JRgob[oHOe4jTH5W7G4ATe;?XN9d<G@gERbQbG0V1[?=^:?aT:d`JFO>
3lHZbZQ3JRgob[oHOe4LHUMk5A0M_M\22Uj9:qg\Mh`U0V47^W3NoMJCX;699bUb
hgCUpj8URLd>Jf_26X>gMqlVblHkfpUMAeAR`;DgmED[V0JaJWOA6;J3B_6V^aId
gc<hhm27p^75K;NU@WoTcBFL8iL70Rn3?YW=<FED;He:LTa6><R?6;lZ[D=qS@Fd
`CdgOna55RN6i40cA`TZGbT`d`ETe:46]AcR_KUQMR47lQodKUn3>Ndh<RK5`[?_
m0dTOna55RN6i40cA`TZGbJ`5\k2T<[dTWJTgIDTqicMBCFIOOLne3KIC_F[>^S_
1RiP>`dQ9\N1nFS[PmWIMd96AXV?ggX_iR5A3DLg0i4DADP2COLne3KIC_F[>^S_
1R5i1=ofoTY6^b2G9EZXZqBSP79AW\Jmd\24]a;\oL8]M?cm1>N\M:e2iCCE6LSN
M<il@@@JFAeWQJ4YIBoS71<YHH7C=ZJmd\24]a;\oL8]M?RCH2Kc7j:\i1CH^=<9
HDp\STDWTYa]l\=G>S2qQ9;60;=d[G=MJTfF?aR8hCj^YO;NC@7Ug7b;:gUeM58X
o@OkcT1U46a>^JGe0;\WQ6TCXA[QP@TZh<AWdd8IPU93@YS5RBjAlJ6A]ddOSEoF
XBXP@8@bcnmGWJGZ0;\WQ6TCXP_iE@>@0o3_]kNBHaAbSReFNlp9V>gDeflFRKXN
6<^3T:lPj9ZfBmjC`Nd<S:jEa80DM63SBj:CO`ZDf:V>ReCf7h]NC<m<5fSFRKXN
6<^3T:lPj9ZfB9n_WAYR\eF86PJ_>KDpQ<<4Vg;@EcdU4MMN3_?A0cGOfjhm<1pK
mn8R;U4[I4OENCXp=1a=IKMq99Rf1HB>QDYFfi`>@OPoe=^p7g`HGBN__2?55bQR
Jh;f2Y`\6kSf8`BMETFgSndX:npXF<_HB;0nl9jk2TM4k=q?V5C7m604_JWM@=`_
HKd;mIngohN_H>d8;RMQgKU1o9Z`d7W5QkSE8UdFg3qD_A:dSN4V@L0GcghUCebD
Jn^ed=TnG[bN0F6GQjONoU_\H1?`9`^g_c83J[4VHKI]YLkSSN:V@L0GcghUCebD
Jn^edcm3kL09bSP:ng0@RHbq[SaJn_j:LK2>gTXICcRbFLWT\>AcaWOS`S8mXaic
70XIPf3W1[DL@9h=4c\J_0RI[>ZV6i69LK2>gTXICcRbFLWT\RFIX8`kU8m]N941
cYWaqX_l^;Tb;80=VmgD:HI524;A48<A<@dPPSAfaGn9G_XWOTJL\TA7KUnT2484
I9MFenl;c20Xe80=VmgD:HI524;O48g@k39>JW\G2kXe@aQfZpS;08TFMmAikNkk
?bP4mlTGh4_fbc5>jM?XSR^lf=9E[OT5Pk\iJScEPIBoE^D;UOI]fYOScdHLYFk7
BQCC:_agPjWZ5541KP=LDI^RH:JQ8E2i^=gKN?j>N]V@eRD3YKSUf[OScdHLYFk7
;QV@:LC_IFnnkAfbY_NRjD`KTqjA_n^>LU7`36mjUAmXXFCA>[>nPT56<XZb211l
Vl_[K8iRA>aHIfai4mYFmSb?hcUEJ`9EL67`36mjUAmXXFCA>[>noT9kk`KlLdA:
]<;UM_pF@AkFUTNhmfGYG;IaAoSCe@F5V;eNJpVX63e=S:?oP1j[T1qMOG1L7mp7
QP38iEiW<S]R\E8HlDqoocYWSn:c`^Nb[Pj7>g?PIadkBDBCJDPOc2pNWOZ84WpN
@jgLQZl_P;<@@j58j\IUKjWkWOZA^7[cBaUCZSO9<J^pG<>l:Gk?Zn4o:TD7i`8a
UaZX>U8O\35YK^i3]7hnbcU[T7eE2_;V2kRM:h;i;3N\G>pJ0`PBME@GlS3c?[V;
N5A1Jg;A;oedT`7MHY]AMn4?JSQN\>l4LNXZ^pESma=>EPZbLA2M2K1jN3B^I1M7
8DXMSjYib5<^GA?H^edC>cb;f81mH;E_d=d70d2j;:AEE<ZbLA2M2K1jN3B^I1M7
Xl@b_i<g\]gQ:mEQ[oq>@B\flJEc<RUB8dohXXhe8F0T9O3NAibLmLZ9>NQb\?9\
e\8gSj1VCPhPh5>eSnj>m>mf5R=c<RUB8dohXXhe8F0T6M_?8K\3dm8\Q@Hh0:Cp
>73AW\=0Pi]b2^NcC1VC1o0A?`Wc2`eCGDPg>ELPDXD`F[cIDQjW?;>Z0?oaVY1[
chLZfCIKPi]b2^NcC1VC1o5c?K:fi4;@o7JV;m4gVkU<qBB5NgKU\lP6@nQ9;6f9
93eN8\9\HH79eOX^F=jiEINc<CBRD\biB4P0h_iKf1DI2BedU0CR8PP:;_PXQ3hX
\I=n0L@<neP96kYeZ^Eo5?K<@0cIKBc141d<K?f3OVDIjBedU0CR8PmNXnPONe4Q
9?<]gNU78o2K1G2pkg8jTL5^X8R6K=_3f^2YVgnQeh9TThB2Rf:6jBUTjMGhXg6M
nEXhgCIZaI<^A3^W=<aeRS5RX8R6K=_3f^2YVgnQeh=2[VCkO^_e0^P\kJlkpQkc
7Ca:4dW0Ofa4X\jT95<TYAWcQUMq54cP0T;2VXT;S;Y1piiC<_d;YdhZV;@MKk^n
o`fnU@J>X[=WBb9FJ@neEcD?D4fkVHMVSe5cXgfDNOZP>E=pioVPW2Tq]Ig@W1]=
E4_PWLMZIQiL<JHK;5QE[Bd1YU=p^6Lh=4Pp;kLA2Gko]Sd:[;:O\JlL7AWpNg;H
9i5a5gb6_L9LNJJho14ilf<WLWJ1kdg]6^\7KZh6poE>aPb7`:;^aUHOMYNeRZ1k
[FfPj1lY50@\M@ccbPVDY8RWgW\[E@hpDADmi_=bodYRF3m?L<5>0<2kWbUU\@KV
15Z7ROEQ=MDU2U0E_ieiDQI1<Yd@D0SbRkGIQl=eodYRF3m?L<5>0<2kWb<^V6:<
9S\\koJU8[c]p;ERR72iOaH5D6SVi>[beNeZYSE5=ZCKg@7=E<U]Pki\a0n67QZ[
HUM8o`J7hS81Z;f`:kfA7aH5D6SVi>[beNeZYS]6?NgR;Ebj?:n>gYMZ;p]dg\LB
dMDnEVCL5ikdl[79LmT2>8^C4^C0?<T0G\f>4D;OgZHVi\1mjU[SgIEg1PK20PWn
SbDnEVCL5ikdl[79CgTE@<WD1Qkn@4jUN>j<j1qK>h@R=Q:^o24nX:Fn?nXCiE^9
dY@fEE@HnOdR_Eh9lCZ\`4ZiL=<0nbDMYmkKGShKSD0SJU[MoD=N2385G8K6cddW
>gm5KEXE1:Ieh2g[H<HTMN9FXBL68k?9Dm62GShKSD0SJU[M`@<n2hM5[\iA61^;
RWgPj:Ch4qHNK2K\TH7JMUoOg`96k:MW=lTg5OE\fK`6h\6[TdBPVALmAOg<WeQm
m\07II2UDd42>`_8TB7JMUoOg`96k:MW=lTgj0W6jdOfS\JH_gJd^kpG8`00MY5;
C@^_@^]=V9G>iBb0B2S@Yq3R>7IFZKZKhXaS=qTIF_He?:`dTDkaWdpJQB_5e=pJ
lKMhi9b:nf62X>2G\I^R1B@oB3M0[j[5A6qM:TAYi[q786nYdTd^bS>6YMi>B[Ei
h:<0JqT=c>I6;MaeL1QQ8e>>]R1ZgfKCP^iZTbCV]PfI`6`ETT>\bGTL1^bPp8Hh
MXZZ=O@d^AdeAgI5IF9>UWU`RYEAEGG7bP^WLUeNlo8nRM_dQnGlZgmdghng];L`
3N_ZoO@d^AdeAgI5IF9>UWUfW__]gG1OJKEf8gM=iqH@LCZ5PF^R:7kSl5]Xd2V2
9DQoQFk7]VVaYJJ\ilkl>YXn=HY1VQU`ldNY5Y<0B6S5MPkEq6Jn44\b65?nHP?L
lbHOKUQcOOA>BPN3<EfD:Q[LKgabA]3Y[[Yi0W3=Y28B25c_]6ML4SYQ45?nHP?L
lbHOKUQcOOem62\JR@6=P<f3@DDA3pOWVVnK<cDZE81R\dBjkSn`X93PE9Pmb9>n
Bl]`VFOHD<FG_WiG8g^QW:QCbQO5I@b?hKdZ6>=ZEk1R\dBjkSn<XOOAST]D==YZ
SY^SKE3LHJp@>jb[?nfb7lIcnl587<8F\G6Uo4P9n_^l@2LS;Ye>NoFPFG8\I0o8
D^O=3CFVjdH@\e]?G^Ok7Fg8IBlCnP=Mm]BWlf8Zb_>[mO;F\m6B`Yg`;PgJ^NG:
54R1iOIDjdR@\e]?G^OkPWhcIb^j5\TXT<XATWO_gUOj<q2bF^]HJa5`9TG8f1Y8
hTch^AS3GNkke@81OcD><?LAfjZN:Xf\4X3[0LGXY5WYENPW5?J7Jf5`9TG8f1Y8
hTch^AS3l>YMiV]j9EPfRmT>E^poJf;A5U[1HLlYbHR]i6?6FF>\5FcUgqVN9d8>
LLUFTG_`>=pOk4did_qdl:Hl<_Dn0F9lhCZ6cHaM@_i@7AU2c^L4A<q__c<mELJ9
V6@ZlRCjibOO<aa79pnWL=MiSq^<d=Fo3F=4C7[<1T7GRmqKH>F\9;7fC1W?9OOi
DKo>6SD@cm1E`F06\_3I>T6M8VmgD5]pPUHW2OjLSA1QK5_?JZbn<;cE>jjQ?_VZ
87VYNLcb35Tm5^AnR>di;_<om9Gl8Q:<eZ0hOOj<SA1QK5_?JZbn<;cE>jjQ?_VZ
5NCJ[EZd=NVf6W`KN^JpHH_b?@DjO?aBKlV55Ohh6P>>BCM[XV3hJ:nl`mG]?L<\
5IoX3>6[4;^3dYS=Ki[XHkH4D@DhO?aBKlV55Ohh6P>>BCM[XV3hEenk7elgI?hQ
FOPnOf<qd59okh:>jVo^N6?iicTb[;<JDiTaUi?UnAP_18cFKAEkj2RVp=fDi5Y\
IG]Lf6QnkekfCCOfN\[@_UEGDIgdIRj\2PP9ocYHSEQ[oA4=3cSe^^=9UE`KBca0
mO4Y3Bk9]FEf<h=]NWFRc5EGo6gbNIO]HSPdGfnmgEa^WiIFjiYPa^9iHqlbmE9]
m_b67TH?VOHiUmZQeF8:0Y@b`3^fAOCL@i:0hQdn8e@kJ;fHb4h0dmEN3DljW;46
S_`gmNbifV1YH>M3Hl8[786L7Jd0gcGE[7V41Ldn8e@kJ;fHb4h0dmEN3DljW;46
KJYg7N_h4Q<`=kMDcKN?p8Wm[W?4h6WHW>K1DJ>naN484g]YRWZidScIX3\KNCUH
c[DBI?nIDTX;[2mV7n`iUjg7m??4j6WHW>K1DJ>naN484g]YRWZidJ_:Z`REmL@j
e9JMB=4@pY;_RJPTHZ28C74UYU4GJC;fM6SdnqaRo5NWQFU>AnDH^\q`08eOX8=l
aS[7X`kfk1cYZ1CqZcC=bmUpHV?;J6Lp`?2QFe[@J2q=NGmDW@K=J`MGUb1IIZ67
A4QUFjY5@05q9`45VKo2Li]IR;Zoo1:GWMn\BcEh@fB75hmI328dAn67m_iH1DJ?
Q8JF]bWFNZSjFABn_Ko2Li]IR;Zoo1:GWMn\BcEh@fB7<f]f\5[`a?@\T@7R<hWq
5lX<IaJUMY^DGX5VOaDU_XV8lE`PEdj=cBeY:Oe\@ihWU9?I4`J[PDiO;cd:J2Af
5D7C4aJUMY^DGX5VOaDU_XV8lE`PEdj=F6eK7KH9cObT6aeN8d>qFo<<ojPmA=f0
G3RR>nKJfeB26c_RgJ345B<VZWjO283d]@[551>e=9=2Zd<Eq=J<\MEMV4S[_g`B
<Kao@L0@`JK=Ad]O=A2kC^m>jfC;UR`AicRCcL`k\MH\5iWcJ4^M\=f_j2]n\h=k
B;Do049ehKdYAYm14NjQ7^J\X[G2XLfiN]6eF1JEUhBX1iAA^qMnchh22keTP281
bWIRf`\h6Km=WHUgRWHBe<PC6LIR\9RMQ:k^cI`4HkXbUa=OOK9CP^;22keTP281
bWIRf`\h6Km=WHUgRWYm];oDIZ1cAnhjA4SP0p@9QiVa@3V0fP_\3EQH[[Mo=Rnb
K9poACiR@mGCBOUa?YkpDKhJ[]Sq37h?L=6pJ;aRFL7q]]ZO9LaqieYW1cVJBKJc
Z^d85n]0AmjH>nEqC^f2j_=q24]Nn]6Y[nKh?hf3k[d3q?ilHZZ=hOLa>U2fH\?i
8Pcd:aneHmc?^<komd3ac@W:m`H<fAaO>R>>L4>IVU[FllL3F`Z=7OLa>U2fH\?i
8Pcd:aneHmc?^<komd3ac@W:m`H<fAaO>R>>L4>IVU[FllL3F`Z=7OLa>U2fH\?i
8Pcd:aneHmc?^<komd3ac@W:m`H<fAaO>R>>L4>IVU[FlcO``7AGbJ]nX2WmXT82
q?j22\PcC]1bf6:;GHBn=I[SmQajQC88G>JncU^mXE^L3?^YfPIT\Nf86bjH2l:H
m?Rf4:Pc]]1bf6:;GHBn=I[Sm1aOLOS5I;SagfGT=E^L3?^YfPIT\Nf86bjH2l:H
m?Rf4:Pc]]1bf6:;GHBn=I[SmQajQC88G>JncU^mXE^L3?^YfPIT\Nf86bjH2l:H
m8]fY:Yh=6lHEJ5;i]lNqIE:HDA;BKaYFgFPLeh\Y93hSNDF8OUa`2l92F?XR\af
K;3dY`k[bG^jV1Z3RXYGoI_L0?A;JL4RF]:nCeZa4L3dSkc83OYMMac91OXXFA7h
Ni2Afm9lEG^jV1Z3RXYGoI_L0?A;JKaYFgFPLeh\Y93hSNDF8OUa`2l92F?XR\af
K;3dY`k[bG^jV1Z3RXYGoN3L8Rna?AjVm6`Pn_D0pBVU`9CIZ^PE1OGZLYjUVWIO
NJ0;_V6aj2kfCA<Ef3KYS<K[]aKV[4M30Ck;Sk=0LI:O:pVfCifZ@;YSRlJ3d@QG
l;eJRX3abdfPWgb=;?020:\aeZNCHe^0TeB8VZRcKePNYIZ@E4UZ@GYSRlJ3d@QG
l;eJRX3abdfPWgb=;?020:\aeZNCHe^0TeB8VZRcKePNYIZ@E4UZ@GYSRlJ3d@QG
l;eJRX3abdfPWgb=;?020:\aeZNCHe^0TeB8VZRcKePNYIIZYc_JFWEV=Y5YZ7_0
Tp>d<OakcW\:`h`n_HONU^KjR=b1Yfpf<PSM\^Tj<ULh5>ep@XiRcL[q1?cil4>i
=L478m08<Jq=NK1`Y4^hPV\:a\QWMR89Tid<JeS1:jc:d6Ffn6TYDHV0WUDq\5MY
PL^lXJCYjH0GE4Y9a4T>FKGO[:nnTX<S>OCMWRCC?02AS3IbWAm3l^^<;CY7`a4[
0L^bXJCYjH0GE4Y9a4T>FKGO[:nn5^X`B;^KBY^GR`4cVYVpR[VmLJaE8j?dO_Sb
5gF^1TOSED>I0@o`adBDJMa?3<:\hdJRKjOfH>]P30jL@9GURRR]dJaE8j?dO_Sb
5gF^1TOSED>I0@o`E3BX0LFI`d8WUAWIMlepnW3a8^2_l?>Lh5EUq`SP_F[[<a5Y
6KcUS3CJ]jdQ@\eaSG^5KhWcX9]Wh:PeDJ]c6I2j=F^BI9F3cc^\JeYKf;LR1[3J
hSXYAb_J2PC40\07c`^5LPWXNIS=YnP^RYlfFl^6``Hjj7?K4ceAJpGM]^kl0EF5
iY^>8@6]hZgWKaYRi42ik<G0agl8Vhn]B:9e86cT9koNA;=Lm@T9\ZGmNU_cmn\P
@PZ[C=@`EL?@c=YnCaFfogkV<G5oRH:hXY9e86cT9koNA;=Lm@T9\ZGmNU_cR92P
@_=@IKOLBiJem@1nqZn5EI1KFT[8NlfBh>:;hWGi`oFeJm82=8\75g8o=8T8@SB>
oXKD4[W>6X2L7EJm?1A6Dd1K1T[8NlfBh>:;hWGi`oFeJm82=c5DO286VHX_2g3i
gjAbpEoQQ;Q@8Pm6cl3Y<:db66k:lmNP6p4Xg070FGHf32`KAOqmhn>kFlp]Q;R0
bmp;Am<`?QB5:ZO5lm[N@=pR15VdHa;P\Ek3e<>7V?m>VGfCl^SDbGBZg\JJ_1A7
hNN\0g^TnTBGmVWJ07P^0fAh_LA@lq2@2f;6E>0[>m:F::O:NplEh>=4DpJRLW3d
V]X@L3oN=4U[QgqT<\=[6FmZ<P0\WYDAdX3YCqX`X:O=0`I]H3eLl8Aon03LVE@i
VK[EOM3JF?ENUe8imQeKREJK_UNl15@^pIORogPoXEMeP\WZjb[FmAn?1d8hogcM
Ok1YH7[9<<WKf5@DA9\[Zd;b9SB\;LJ3Y:gO_BPohEMeP\WZjb[FmAn?1d8hogcM
Ok1YH7[9<<WKf5@DA9\[Zd;b9SB\;LJ3Y:gO_BPohEMeP\WZjb[FmAn?1d8hogcM
Ok1YH7[9<<WKf5@DA9\[Zd;b9SB\;LJ3YP2WW]7bgHlIViUS<T2>p1okVTUHX[CI
DjMQGlXC[_R>NTSUQc^EJJW?@:nP:WYNbOnbV]ll;3c?e2c:Iib]E1d6hgJHl[CI
DjMQGlXC[_R>NTQUQRB^LNYbiJ9b<aYN=OnbV]ll;3c?e2c:Iib]E1d6hgJHl[CI
DjMQGlXC[_R>NTSUQc^EJJW?@:nP:WYNbOnbV]ll;3c?e2c:Iib]E12\\gX\Lneh
FbAZQlA41phajJNc7KBCZb006Z]do;@7YYe]X_SGVESlLkd]YX43NZkCeLnTVEL3
5b2<n_O2OSho9kT\77BCZb00R[e]Kj@8Y?8NOCcGMEL@IDd4V24M3lJLa_0IlDC3
5b2<n_O2OSho9kT\77BCZb006Z]do;@7YYe]X_SGVESlLkd]YX43NZkCeLnTVEL3
5b2<n_O2OShYnnT[H5DcomaSFRFLmiq[11W8hD[Yc?>MceaU2l;@d77E[R49D:2X
2i6Uh]d:SK:[nR1iR5\>NM^I;dgkH[YD2l_U1DgYc?>MceaU2l;@d77E[R49D:2X
2i6Uh]d:SK:[nR1iR5\>NM^I;dgkH[YD2l_U1DgYc?>MceaU2l;@d77E[R49D:2X
2i6Uh]d:SK:[nR1iR5\>NM^I;dgkH[YDWo_fVlVfO^8gPm1MRklpGON@`P?8_@nL
fmhW8^_9U0nK\1H3[[pPBZ;AE0SL3M4=SJ]>[qf`XMV9mp@Zjn<^gpGF[_lg\4f=
^@WOB^[e=bjA\qZ>J>kP[JTHd>145G9?UNQa[G7BTAR8DfkfFc^YmoQ?7`i[mRX[
SI7]HecgcbY`q=7cchE]Va]`N5DEZo8`gIjE8Dd[5ke4Oei[eVlJ^L52H5i^FF23
[GVX8jg<dJ:6cYX`<`E]Oa]`N5DEZo8`gIjE8Dd[5ke4Oei[eVlJ^L52H5i^FF23
[GVX8jg<dJ:6cYX`<`E]Oa]`N5DEZo8`gIjE8Dd[5ke4Oei[eVlJ^L52H5i^FF23
[GVX8jg<dJ:6cV9?N0R9g[ofmgDSTQX\pSIgSZiXKFaXWe<J_1PknIiX``Y:<?eI
XBJ^CV\M@`=8<U_0:fCgfYDJn8De\m<iIS5CEV_XKFaXWe<J_1PknIiX``h:=][T
Z2n7BkDbd4=8jU_0:fCgfYDJn8De\m<iIS5CEV_XKFaXWe<J_1PknIiX``Y:<?eI
XBJ^CV\M@`=8<U_0:fCgfYDJn8De\m<iISPDSVR6o9AN@FC7i1:;_p8j8k^C:XCN
Y?3SaV^MX]a\>[`XkNCT1PPGV^?bMTXj6G=k5b;RW3WV5b9eXh2O4:8k42bcL\1W
Y8D:a`^MX]6KkC;hTQC1mnP[@Ua=MZj7joMkIECRhF<ZiKDb;W8d4l8k42bcL\1W
Y8D:a`^MX]a\>[`XkNCT1PPGV^?bMTXj6G=k5b;RW3WV5b9eXh2O4:8k42bcL\1W
H5O:@\m@?]6g9d>IXIT9qUm97_X]E_e46_k7JJDXWeOJ=l]]GXO;EWf?ZhGcO?aH
^\cjSnPOYlnB0el59BC]h8T:\e?]E_e46_k7JJDXWeOJ=l]]GXO;EWf?ZhGcO?aH
^\cjSnPOYlnB0el59BC]h8T:\e?]E_e46_k7JJDXWeOJ=l]]GXO;EWf?ZhGcO?aH
^\cjSnPOYlnB0el59BC]h8o^91eFNcOd8G>6L5OQXp<Q3Jh6AcB>FSH4W>eDY9M2
1?BHmCSKpeYB9gX]K2R@hPZT;kSp4IGQ6L8q`ZS2969HYL?4cSnNb@DM=ORHKI]]
<kblkBNa3<LMR55jene?O3^@h_MRjBhAP8NC4OFlo=@=3i=Kj342>43QQghShWgN
Zm5WaOVh3Ca@15J@G6D>YK^FX<f[90h`Fk;\I3nRn5D>nA?=1[cqR5``DfC5D;[S
LF;eV4cL\AL=A`QYY?3SiomiEZ2OEd1>8GMWETC7RX1qm7ocSOh7`N>dJe=H\;dO
T5MMqWj>_R>[?e4LGh2F9OHC\\9:mCYD6V@]b=;Aoq=3WTK0SHp1J;oNIB>0ECdY
YIKg6fCQYC6VEmTVGpYH8hFmaYAo1TdbhVaL1j^JRo8MWUn?k^I72gHfFnlZYa]Z
BPfV?JW;M?HLAHhCOeJ0cEG>aMAo1TdbhVaL1j^JRo8MWUn?k^IY>Emk:m6ch3\Z
B4fV?JW;M?HLAHhCOeJ0cEG>aMAo1TdbhVaL1j^JRo8MWUn?k^IY>E3i_\h=5gAP
jAH=?Mp=SREg>HXUo:g11Tb2lN5c@@=cWF3:T<8lEmLe[KGVS]joSH@eXDClH:Lm
^p[<5Lb061U3fWSQ_8J0of=H=LDHg>2WWj;G\[0fXD\KMKBH5O\n9B<\G<KR>=@O
EFXXhh766@U3fWSQ_8J0of=H=LD4[9hNa^?L;BRK_;`inG59FOcf9;<\G<KR>=@O
EFXXhh766@U3fWSQ_8J0of=H=LD4[9hNa^?L;BcFoo_IDONdo>lCImq0cZCB>daI
5]jbIK3`f4642f[<4UZoTekOG8R@h6k9JlZ_dCdkZ`b^3iOYmo:\GmnoE:i7gdOI
5]jbIK3`f4642k<ANa>i1X\@fDFMO6CJhWQbZ_^e]G`A9ijYmo:\GmnoE:i7gdOI
5]jbIK3`f4642k<ANa>i1X\@fDFCUZ9J1c<<_gm<cmTqMIAGK7mSVDeI@<=LidQ:
BA[e96Bollg88lC4bQ^\]An06d<`3nmh<0PgAfdDJ]7a;_j?FlmSVDeI@<=LidVo
`mfHS9LiL2a]XARIPA5eJ@9;NmdQOGG_;1>6AfdDJ]7a;_j?FlmSVDeI@<=LidVo
`mfHS9LiL2a]XARI\V3k4?<N1EnG?iE[p@_MQnnndCX`M7bMGVAYQUg<K6a0PQh8
EDJ702QN2:]aWM7H_?g9]bnA=1M>T?];AH>]b0an7CX`M7bMGOY_gOSYF;GF=D?M
bS:Sc_d;k`=\;Ye4fm\?kXbST1M>T?];AH>]b0an7CX`M7bMGOY_gOSYF;GF=D?M
bS:Sc\;RXYaoX4Ye06bRgp:3];62`M>]4JanYF2=^]0AlI1HBSg<Zda0CWh8_WJ7
a`QNR5]amE7H2b\?m=bS@NM>A2]91Wg5b8FoLhBbk5Wof9Y_ORSYjXGF=S?MRG:S
mDd;GL=\oOe4oc\?m=bS@NM>A2b91WC0m6anYFX`oJbMfMY_ORSYjXGF=S^AJl;;
4RHFP:\74>pP\>1k;5=C8Xk7K`j8<XePAWHH2_<mHlJ]0iCTA^5f7<1fUClX3bOQ
QbZf\C`cQH2PU;LBNo`O]bb1[e^8<XePAWHH2_<7MUdL^^dBD8XjjeI<AUA`COk;
CWodDniG^bEhU;YBNo`O]bb1[I1fb@o=Z6RfC67eCQa?R7i<\TAgdFff@73gC5Bq
G^h_;9K=ScfUUB5i41`6n8B`kJBJHbSR0dX7N3B^jWRM6S<ZgmkCif6^BUaoDI2T
GTM0LKZ4^PQ?5[PCD]SoaJBXkJBJHbSR0dX7NT2=JbJCLBNk8TFT@<^;dE49jI2Z
GTM0L2cnLgFM^Die41`6n_E`4j:1_OgP=L@GVa[i?OWX0T?2@5?PpM:@lKI<UVL;
V`h_YoSbKq?l2dkQLASokBK0i:1m>UC>]iX@K;d@d;i\^?Z]8US5jlB<\[b@14;>
0bfZf`[fJHFmX4TdL<SokBK?YA0QJN\_MTciYOS>6ik8^dZ]8US5jlBG6c64Gn>C
X^:ENnHomV?Pn^]nTBf]1lB`JI1m>UC>]i4YYj5LBOZjX3`I5;am2cH5>jL3l?pK
a8[<kj=bgCbZn_V<V_EGKlBhIE9DmcU1f:j9K@a2UUDl]HoaFf7YW?V:KDkGXQck
gc[3@j6bgCbZnJ3KgPa8\^;:eUJ5728=na6AaTFAoUTl]Hoahn5JW?L[eJ?E75IK
<4Y1MMTGlG;mDO_<V_EGKlBhI755728=na6nOS<7g:?TRY\?LJ8pE^F0nei^OPaP
8GO49=YZje>\Vc4Ab`TgOl5b0h_LkoTjH8C\:i;EAnR7fkK6XJTg;U:ghJiQOPaP
8GIE4P<MAKjSS]1L7X=dSeJ2=_PdL\?b]8XhI=UOT?3C4l:an62_E@Q3jZ?TTQ?1
E<5d9=YZje>\Vc4AmX=eSeJ2V>M>Pi=J=>Z[oHgSpZGkLBB\?>RWSB7;nIi?Kj=G
86_h@cB^G2FjigM8jeCaFV0GNZ1M483o06Gmndc\Pg9^GVb\A3RW=B7;nLZd`N^@
jWAnYK_;0Q1hXl9I<?Td432\E7gmD83o06GmnSk2FZJ7h]RToE<A`amSjXi?Hj=G
86_h@cN;4Q1hXalm=NMiQ;@[@f_3aqFN_Km`SFFY7CgU@nhc6M=0i_eeAJP5UiEa
adlK2fW760`Ea84h;430XGlL1dTbnVF2nIT3SVFY7CgU@nh2]KM0WFCS4KX9Q5n1
;8nm6L@A6fk1>b?CZkL2X@lL1dTDkYFhiEdRkB?CP]V5ZdRJ;U=0i_eeAJPLPSn1
;8;XJ[YXiClZ<YjUJOpYi6[CIKJF==kiVBc^2O[1a\o85nn2f3\ZPmgo6de2820Q
?;LoT0]c1jm^mMeWog5BMQ<k@KbF==kiVBc^2O[1WOYSQO=mAVWaPmF9_[7CMHHe
LIndKY>A827H=MdWE\5Y`76?ZQA^BH=K\SEODMeXj\A85nn2fP\cEa8^NRfli0LL
7Um60dbpTf>PT2Ic4P<MAKjSS]1L7X_H8l5l0h_L:k?Hk8XMI=UOT0=IEl:_n62_
E@Q3jPiAOPaP8GIE4P<MAKjSS]1L7X=dSeJ2:h_GkoTjHTX\I=UOZ=RTfkK6XJTg
;U3ZaZ?cTQ?1E<5d9=YZje>\Vc4Ab`TgOl5b0hUQc\U;Q<7mK3LngdSFfef_q0]c
a_>`U7WYMbH6iY?=q8GNdV_FD\]MJo1_5jZ2^M<G3Pl`@OhIIFB<EaOf5AG@@Dh<
>o@<n\b_ljM[e_=BeLUeb:TFb\]MJo14RjZ2^M<fLfUUJR69kNH]BgOf<AG@@D48
?b^a`726g>iV@GB>T8VkQo3^ihf7gfK7BZhbh[NaCJl`dO6QkbB<FG0?K2ZngX0J
A;ZnQp>Y_K8@I\[_oO7giOaYkgfWkH<oEM?BZgL>=TIe`o0X6ZZ7Ha<]@_gKFF;g
PjXC:NiU\[^iIXX_o[7giOaYkgfgNXO9Mne^7^NZe=Ie`o0X6ZZ7Ha7Lk0YbiP7_
h8;_:XQI><GTjC^Df5dmfbRHiG5\kO<oEMe^S^L>SGoG5C:3l3igHS6De0q6hGNR
IJie`N4_J<ah2gn3[l8NPU8Nkn4]QmOLcCj`??b\?W6e5lgEK\L\lUM]D]Rml?Qj
WJfe`N4_J<ah2gn=jdYUlUQOlWKAol;LcCj`??b\?W6e5HE6<RQRd0c]D]Rm53WC
Ha946JU\jdR3eP4mdlkNPL8Oani]Q>Omn?FQ68b<ZIRnQf2p@[BBfoFngN`UaTnN
hGCIAUU`Ei03jDa`@Vc9g?Fi5iNTNI3ahA4h;Ej=`]7IJ<ZEBSER`\F2gN`UaTnN
hG3ILmR\iiVG4Um8RYBGcPF85iNTNI3ahA4hZ[knL]7;J<ZEBS``j@l25MdV\f4[
kO?`AUU`LkPBjDa`@Vc9:E`ZB]\o=>R9A7Ncqle[]gkbBHIY>@kejGh>aUn8_6Z8
2h<FE1I\21?iZf82oPENfcjTOL^oCE@:=0YLb?K@l57LK\fYX@kejYZT>O3L<6ZB
<^`XbUf]44cQZ582oPENfcjTOPQ^jE@:=0YLb?K@lo7027XmNXU_7:>>aUndPWB8
Uh<FE1I\20X[]<_>OA0d9hAA4p0^IK?]MO1FVBU[bnPi]b2^G`3[o:mK9aAL@AoR
Ngo[H9lEFLm8U^YOZ5PDedh2>`OM>iJ5D<>?LALi<On4W2HMC53[o:Yo5c?_OhCP
ElGoLhDEF<mPB:kOZ3PDedh2>`74@YWJPi>?LALi^OPi]bQ3Ca3[o:mK9aAL@Ad7
H4nfEh@_^_2K_Lq78[8kdI3cVPc3KJRLjA>7WiU_5Cmn1@AicUReIIZlnAMi_@[W
ioHEXF^KNY4VW>XIQhg44U=`:nEj0JMLjA>7GOK_5CmnFMaK>7<8[LPZdSZKal@N
:c=4XF^KNY4VW>X;`[;oLd=`:nEj@nH96i:YWi[_5Cmn1@AicUR0kLX9=3OSCh6e
X=Opfe<HPZn0T1aRo8ZG@Yfgbbl>:eQMYNNZXSl>LZA2Hg06XIhoGQ=JB`WNEk:E
VH2a2kIih0J:p;ecMcC?cF]2FRlUebDi_7YdXNNhOm\=VLY\KfAL\=ZhgKTU>W_]
No8aSTUK[0ii@BTGhdW@e1E:M4MU5bDi_91e99Nhbm\0<_eG]<EF?^1>neL7_J@A
7o8aSTUK[0ii@B3jc5\?h4E:<4M1\3^oO7YdX9Nhbm\=VLY\KL^l_dYe5JOeMKCB
Rq1bWFT==:YX1LQL6S;CkOM2]hikEm80]bSJD=lfbh:8NP:T<Dajj2=dfRgjU>WU
`X]fJNL5J[`bJEWL6S;CCdM2]h[kEb80]bSJ4EC>QEbg6<4hFPajj2=dfRgjU>WU
`X]fJNBM=dYfJ^WLHX^8kAM2]h[kEb80]bSJD=8J@c=C\48:kA;W8?q@ZY5O4d:D
h:HJJ;RD\jGfB0;C^JY:Xo5nDif_]0OjRm]Pc<UJoV7hHV]g:\3ATXTl=Ck2]Z9o
<D3JJA7WejffB0;C^JY:Xo5nDif_]0OjRm]Pc<UJoV7hHV]g:\3ATXTl=Ck2QdCD
n]NJJ372\jDfB0;C^JY:Xo5nDif5jg^J`H4@dUU48imqTAF`06^Llh96W1P[K]VW
en\XYFT3S^J5RR2DCJFDGa>7?gJ?3h7CgPJXmb;E7<D\cd3`b8mf`0NV@A1a>nA\
4n\P9aDBBenlNOEkej:]3k;\Pf2fiN_9Sl0Bc333lV6Ed5YnUI^ZlhPC@A1a>nA\
4n\P9aDBBenlNOEkej:]3kRO7mCl2Y7AWl0dc333lV6Ed5YnUI3]ckIKMMg:jh0\
=<1pBdFMY;C:]8BTbNP>^;?XchLYb70=ej[U>9Sq1dT2JIaRL:\fVl8^kf0\:ZM;
aTJhoVWb<Q\ON_[`Wd<<l:@6E4iLfjJlRl;gP@R`iDMfESlP=?:oblg0Qf0E:X^Y
onH3W9_VmQJnKSA?]TC8^KaQkE4Khj2VC[l:`]R0Ce\F`3aeL:\eU6GmQf0E:X^Y
onH3W9_VmW^m6GAc]U5KQZc^=dK1Tj2fC[l:`]R0Ce\F`3RoBRcL^mJ9KRSBXALq
5<0_QMVg^Di[E2ZJGZKn]@L6`aNK>_PV_?2YG0IF^7UCb@W9j>]eGAcSn>c]E@QF
FoY_9g6Mg0QeooV[GZ]no0cP_6jeUWjjBA`T36Q;^Uo7ZSJR[UO2CAhRZXLX9g;?
fT6M_CVX^C<o?lfJ\GK6YSck_6jeUWjjBeFGDHi]XN@d`1_GV3Vg=kaDZXLX9g;?
fT6M_CRX79R9A7mL0k[g`Rlp3[kEmVjEZJl6^5_lV46\e03dL^X@`Th;_;n[ckS]
>aOg?7W:fTMLOTFi?OAhMKc8O4]6:Wf35P\^QjC<fLnf7h^6CM\MOPXc0[Hj7D][
1fEGb^;XF^jYL?79m\7JEMj6H3CFGjj74Wbf`j<497RWU03N9^dDKePQl[j^3kST
>aOg?c`^9OPoZ6KkNKA<5Hl4O4]6:Wf35j\4QjC<f8J?7h^6CM\MOPXc0EQE7D][
kY74[cBKmKfKDVncm\6OU6J_O[C_kk[d;ebqC>W5bP^h8bMaXjlh?7lT4f?:Rd7K
@K`U;KjTSNf>h7l\B:eF^6<7g5Ho<P;8PSgN@3ZY11[dkSdh3\ij;KI]VT1@ObRF
O\>Ehm438k42bcL\1WY8D:a`^5QS@`40?HK?TiKZXJfZ62A>]3b71?@8kf=XnEEP
V=I2PIcGSNf>h7l\BAm\RnCMeQPLL:84mmd8IU\mX4^G8nV4f[dCNLG2;RHcMbR4
O\>EhCg0d4ZAH^_e`Z=`hm9OlgJ:C7qOW;2Sc:QPa<2:Lag>J0k0IJ_D[Fb<?KRV
hGWnYlJLGTCUEVXAEmSLhCf3iiN\linN3Gl^cidBoY?I6\ZK?8FjL3:Jh<=i51F1
>CdTe^2hDKYWSL58KU`oU42B;S82LU8H]32NebCLoYICRAYDNMgmb[:k:d_<ZGMo
L_hnYlJLGTCUEVXAHZ6K@Lo?NDV^Oh4BQ@la=:YPUGg0FMNFA8<TGb:gh<li51F1
GJ@=FBR8TU2jg]]:c>mLg=`7QqJgj;<dIf1YJi9l;U\D`n2`DNbZG6Ph1a7S_>QM
`M3D_9Gi^527dB[?omZb6?`OCmZ17feJA<6OO\fI@TI:;C:ldJnO==^dS]>eSU\E
A5eAGiPVZ>\C`d6GPeOS?iZhIInNmWnNLE3Yo;g50GfL8J6Cf@f`l:bD;>5eVdQM
`M3D_9Gi^527dBDI;jXeJYb2<WfhlMZcIZ1TeXeFh^\\lj5LDD5O=N^dS]>Tf5gV
VMhg;iTFZ=ZF<WmQ9hXJp^lbiN8R<ClX9VX=@9GEcU:Q4YI_imo3neGGk2fb0E=L
k7;cCk_JH7afN2mo_j6l3K>jf3<Tgf8_7A63IMfSB@X36NbA7An[JB7f^B;h@lWU
Oj2b@]1L>>hNUM<i3VoCXbEP1E5>7:0O;Gm]`V1MZi8SBXdJJHTk7@FMelfbAE=L
k7;cCk_JH7[bM5RJoEgOXVQj65;e=C^]OoOT=9GW6OfSgPbAPAn[JB3F7EZn5ZcG
_UfCI_Kj0lD_JdMp44GQ6EQLViKJ96@Ua6cW5F6e@EoUDNWekKPZKbF74bl[VjRf
^XXeKW?dj@m>2FGB6L1:cDNl2EHCGn\246c@[T=R<AU_UdIBTTha3Q;?b6<MSQRT
n3f801\mf^PB<IL0Yiio1T=6b2bTG384?58M9I1H9G^UD5;MJ_iZbO9c4bl[VjRf
^XXeKGWe4gjD=1H7LGIdF8]1biLZa>f=a0o;YZhO<AU_UdIBTTWCQTSPCiToX[5Q
06h6ToHOHYpXUPjU:O4fP@l7N0>`LLdg2N_9]0g\4M;8MD8_n<`Zc?klbiR;R[E`
2PPVaPHSmlPGV:<R3SpQH^4fHT;_;HbX0a7<;]oOSgR5BF16hZl:PNOh3DK=<iP@
<SRTB0h7JbX@GS=dZL`JoO_TZG1Q>IQA;lF@;]COSMh:X[8Z:Ikh7]_K5kh>QMZ3
3D4;B6;Pg`XNf<ckUM`F=>I_kMD\:CX9N]Q`Thkj2DS7MN:oZZKQ\[_[m94H<i7@
<SRTB0h7MjXIA8`PQc59N@Kd>a4CkgIDTlm<g9=5E>_:X[8Z:Ikh7]_KWe6@BAFO
<bC9P]gZ;DGg9p>f_h_?MSd`2V8HSc9oA9;EmBG5hjef]I`ha@:`m6Yi4J;h2>;=
hIMZiLd\nEjf0X4CTD=DR^>j`94hKX3oA9;EmBXieT5GXG_LL2n074eBmiahnXb=
3YemO@02KOS=:27YNZX]3GWKjWnWLE6<CFh_i\c@OanFmJ:1n\c3^1enZ09Q2U;=
hIMDaL4@D:;ATlL:TfUG>Sd`KhjhKE3gO>XQFFXieT5GXG_LL2n074@O6hQLHZF5
Z0H47ciaqCEHD[M3A4D]9EFn`iM1E:=9A94NAfC;bXhdbd8I3eIRRGPGh6JO9?;]
JMYjL@HCJ?2Fo@WMFSdLfdFnki]IE?R]ndOjl4CBbIgD6bbold=SNV]@52=YGJ@a
kh?=47mC>o5;b_n:]]he5@VeJclk62S2bXZF=mm4boYm2d8I3eIRRGHWK8MT`g;]
JMYjL91kTZnho5S?c[=ZcY>JnDQGHSVWq\c8nDEBBQ2Ke>lm9m_>dIOB;]O=PQ^D
YESG<M2:e5glj7j[c_if1N1NK0Nh@Mf37\mfJ\d;mKU0@ACnoZ;[EQ]4@fY@RV5D
V[Ug^N:KNd2AMFOkVh3`Sb^U@0THWiI?jS9A?BkheW70MAlPBNl_fQ`l[LF_YjXM
;llbbM2:e5glj7Ak8Z[`2NOBiFmVC1nLV3^PdnZP?clHE3J1X9kSV\=dqfZC:]h:
Hifk2C<8LI[JCi3fJCEB1NPI`h6Qbi:iPKXH1<j[7mKc@A0^8;04JFdC[PR\eTo:
Rifk2C73<?S==C2fR[EloVSf^hBIaKBWDR>Do?3Q@SDnoaAG0]KY9L58YZY?2Co^
OlS<9[;5F]iNSPYARKd3Q@JLKDBQ=i:iPKXEon]5omVP4Kl^_j`6NgI5>nR\SToO
mgKhNUWTgXNh7<0nqbUlL8;[;>_mWEi1@85GY\VE:fmH<_LGmo>ZD=?66aYNiWo8
k\;IkfhCni87RFHgg9M_MGI[C>_mWEiD<hMmN6:E6f4375c<_o>ZDbgCjb_3Lh40
?`I9^2@BiJJleOS3?gY>1OV?YAlfFOIb\^H1V`[T3kN9cKXAOo>ZD=\6b[\MYmo8
J\QCc_6O_n:07FHgg9M_MGIMjENgT_Bag=f:bKSEqfZ7DDef>[lCmKK:FJ5]Skok
JKVj;D^P?>KJF\lVdF\B]^e3?VklNNL2_AEDTQKU@]f8ZZMfb[lCmKK:FgYnSKD_
PUmQQndRd>KJFOeFm?kJ02A\DDRC]1Uo791Cb4ZVB23=GdmjD<0_EIO4EiHI4EEf
UeS0U^^PZ>KJFOehJ:KDK^e>YQkloNL2_AEDTQKU@]f8ZZM1G^TbA[CE6H4KCFG]
p=bnUFH2dn]jZjCH[blNUEOfOLV1cU4\T5Vb4IO]Hd_UkVh6>6Wo>AB2dW4JLgR\
g;O<6=l2dn]jZjCH[blhUa6fk\[@_F=\K<3Y6N\j8SPUmVh6>6Wo>AB2dW4JLgR\
g;O<6=lLD9[a7BSH_blfUC6`_Y1EjU4\T<3Y6\Hl:=gcKgc4E_<>Ip=Q<SgT_iZ^
h4:NEBQULjX74KCQa0cJ5fN;C88e9pUTM`YKUK3l`;bjH[\03<E_10>O?=kI@3LT
GLoFZ8P:TmUd5e[:P3fbho\O7^nRWc`c14<hUG3VXEhWQ1SFC8dZ1K>OC=KCo0S1
oXc1`YP:TmUd5e[:P3fbho\O7^nRWc`c14lLL]AYPDnjHF\03<R\mXSjAdSCoQS1
oXYXO>VX7fTM@KlP\Mq4:\;5FHNI<;PV[HlCJLVU9nfh;dnI3>?3iF@B`Jj]Wa3K
_31Bn`e\2QjHOnheJ\W0Jghc1CCm?@3Af^TUjYPmY[9HA:SW\JLih:Lo9REAaIHJ
A?>a[TJoHf2SLV`;;b60Jgh?2HeI<;PV[HlCJLVU9QAkNCeKHD]VTK]j@W2W5;bf
_31Bn`e\2QjHOnheJ\W0Jgh?2cX;GUASZ1O[_:jgF1pH1VEeC3a5^i]VD>:8l;gK
HT5m1^17eR2=]e_m89;\3l778diMR?Ymhc@Lh7Ll9Ya:VTb4i3JEga7cOER473fc
X<`7M`9hMGa<>g<Ih7=2ZTP4cIEl0RllhkU6ZQ[C[2d:`=W;_3U5^i]VD>:8l;gK
HT5m1_mjQlV`>64IL6;=LlN78diMR?Ymhc@Lh7Ll9Ya:`=W;_QNO\mhS3b7NaFE:
Z0qe3^j^1N>`bog;c8jg_ifRmUKX=2PCKTZJV=@oO6]ki_>0QSBXGCVYMMRjV[i3
0R1^M8kaR3:]=72hUn6k<TVURS7X;RCC8^ReL@;:dGYA3ffYI`]c=QlFePKh89bU
8ZR_=8GIdNM`bog;c8jg_ifRmUKX=2PC8UZGV=Do<P7Ai_UF5iXljCZYMMRjV[i3
0R1^=8OIdSMH[kNP9ak9cmYDIXq;`S8m6oa=XSM7Z\L\GCKTKCq:bN[dBXmc;5oA
H9\=XTSmD>=WS=F9AM@bCh?XKdjX8H\o<?o:XQk>O@e^5GYS_L]4ObgfoBB]TKP\
:fXU\KC748<2ZLfJ72I4CJSF\KG[X:cT6]BAfjk=ZP1PT690XfVbn06C@X2c;5oA
H9\=XTSmD>=WSLB:>750K6KXKdj]jhgY3oHb;EM=XiO^5GYS_L]4n0eC@O2oQLi\
F5>?H4hH56p]mg[OJAH@T`KOF6C5fV5JH6:\KOdahjj`]O^Pi2`B2m]o>3eZnbaX
aP<iZD^>;]d>MU5^D0Y0oF<dbWNO8?\E;[0k<R_ahjj`]O^[>m8F2W9Y<]_HA[@=
U1_RZN>1Ne;kbW\<UNVh<jk8AZ[Om?QMb;N;IFJ@2W:ho`M2SI]3bn4aTO7^kV;j
nk=W7@:g:DK]cN=XOCBJ9`BOF6C5fV5JH6:\KOdahjj`]O^[SI]3_SfB?`n;_J`D
:@CFJqjX1^3F6[50PeM;b58?ZdIMRO=]?\RQ6eoJQfC?FJ7oS>7RITG64KlF@[W=
WgclXX`0b6GMM2:6HKOf]P:8>hfb7T>cPeIm6FoJQfC7]Kj:FCY=<L2o4:lJRb^5
PP;l]3E6\0X:@7gPHDO]iI4MmOIMRO=?XAao@jCL^fCWMklXnVfCPX`6Q?^FJiF5
<NcKBW:`JMIE`5Z5gBAIFJCDgS56TR>cPeY:Fi^nO:lEKZj:>kIYCILC?2FGEAH=
7[g:Nb2?:^gS6750PeQjlR3oN6fK>oXF?EpL_7CAfI8ofi3WdAAJF>f\cSQ4l[hb
iC45i6G_6Dd>?_gH^UYH\QMRCe@VanJWVa1idEXRWKgp:Y89c9o>h1IXh:Tk@[@C
B1APf>\On7I6Y^[6T[LR`C_Bn1YAnIdd[m\g>?nM1VSRP^P1[WdcKoNJT:\>kaIP
YB8a7dN;NoILY^[6T2W2>8d=9^a_4R;7P\l0F?1ajRT\O7j6nK8`3H9k888YOanh
B1APf>l<hOUo>?oaneeT>GIjDeQ?n?dd[m\g>?nM1VSRP=LTOl_mAIRi:m=485YS
G2_b2G^3i;lE[;eilZSj>8>D^YG`5MNe>acF_Q[k[9\Hg8K3@\ojh1IX36<>m^Yd
JY8S=Rc@qFf?89Phehj92JGc>NcmgUcT57D\:?fV\LomRNT=cJAUO1K=4G:dUh1c
G4ZLWnd15<FmDgn<Za6XJS\3Sck@Z5O\f<JUBdHPo;SKii5aKKgQiVT4Mk?A4[QA
=9mYdK1N8`Q1JEQ_n>ehj2b2?mW@P_cT57D9:KfX5J=YoWlVOOB0K76U6>H^JQiV
Vjm9NcdmZjT1bTBK[[<Je>7RSQUVVBcTA7D\:XHEo]anm1JaXKZh@0Y[]Ei^Xl[3
JLUN8S`KAZH`Mjkhfhj926;b>LbI[F>1UUME@p=W[?3gPC?P]GJgBPlX3JIG@T1>
FM4\D8@WM`Q5Vc0;2TZm8@Z1DL6AOB]5B]J4[Zm;Vj?MCV3=6o7`:XbFHnIMi[P;
PNN^H;d`?<_D_k5BB6K^;\iP3Y6VOBfR4Oa?DnjLQ3ZDN3=_Dj0Z16f>Oh4UifP5
S7]?[6_L7JS[Vk0;eHAJjMiP8e8PkCIKBYT?^mjaX406DNV`h?Z`3nbBJnbnL16J
mkN^H;d`?<_D_k80c4dm8WZSH1k@dXmRDCDW1E>`9DPCP^?P]GJgBPlX3JIG@T1>
FM43=G\3K2:i17m=Wo4dp4L3NUUB<H6=AKOKchjI?]O7TSIG;bnmSTO0>kVZ=nfF
d=mjZH^2kEI2bAa1i_c=O4l8VkX9onZ^h@E@31>6Q`B2M>^Ta>>go2MM7\b]Y6E0
`bVjQ;^>VIJGLTA6o\WC9<N:EDBfih;ASYFcOW`7X>PVbOd5J6eaF>3MX4cOLhPW
ClHbX:D<^cNZZOCmj^h5J4l8VPW9UH6=AKOKchjI?]O7TSIG;bnmSTO0>kVZ=nfj
`=AJM_Qc:HVk46WMq<T<>cZLHMR>=SmbS;G>:\oPV4oc:?me0S@J=>AR@;`PF]m6
^ceI[e0]l6U:Wlnjoe6^VWEVJHSLI1icNMQO5IGIWEK3H3WFDHAhZRbY4Lcf?D2`
mAk];`oINM[_SbBeATkCW8<5BT[L^]JNmQQWa^]@i]>jC<G]FAm6U]DM6?[4<832
bceR[=^PJAlmMHBkW<iN?F=LFMR>=SmbS;G>:\oPV4oc:?me0S@J=>AR@;hZfaaV
c7nUce`W6@gpGA6I62?9c]Zl>9mI]@QEa^iX[:ZoBiJ6H=Q[J?1\84U_R\;6164Y
ScM`j95jaon2Rai`KI0`akHQLF44NobAQ?GB9XTj^1NeUC=[j1k2moFDAA<5Cm]<
H8jn;L=]5jTNYY54Y^7dKXhcLbC;_UEP7jQdZ=ePGXO6lB[=nm>?W51>i>n0164Y
MD1abVE=[8TLCD34cI?dc]Zl>9mI]@QEa^iX[:ZoBiJ6H=Q[J?1\83nkeW6Y3lb?
WNh=ADpG?G\lFO<=TVRL41HD4PecfTJOUKAPXQMICaXhBB`QF]lI<4KT92;7C7G=
>5ma[^Afl=O>ODS9Z`S[4fmKcVGOWSj8aPA9Ni>Aha:YhXHD5hnNj4lE>FoSFR\R
SH_ZhkbWa1Vbj1<PGbab47cZg__BY\nY4=Jm06Ajbh1V6l\]>1^EAn=192U7?P\a
1IbJ4BI:_^]QdOH=TVRL41HD4PecfTJOUKAPXQMICaXhBB`QoU9b6[1^alYe?NK@
9q?BEGC3`N<bZh<M\3U3eDIG00dM`QSSP4FlAjJSm_CWMhANAXOHA]78qbHTbhQR
TY:;TBP]oM<4\l6;5Se^:LL0nHoMh_PUkGW6I4h]U2T=Z[OV>\VK1V0Z`Z;Si?04
L5XA@@X]GE3bkb2N_R`VT:S5fOWNhVfHXnndhS27HS]iVYTXfEYDEUe6PE9Qgn6Q
MiW;7oX]@EgI;nakkkQVJXn^F\449lOnl]I;4TAmN;iUKafXVEYDE`Pi;X:nY;^R
jY:;TBP]oM<4\l6;5Se^:LL0nHoMh_PUkG1l9Oa5W987`MQ06YhpmeL\>MFoO;jm
_X6gaZd@MP3LmLjomWd<^6N]FSA:Jc@m:3MU_e3N82DbMWUh`>@hd9M`E[5?H9Ca
gce[kZhC=<f[FF7C><nWUhFVH];O`8jHjoC05@V7FPZPeM?eQh8EQ>biL[>bPX8P
Aceak;W[7Rl@`b5kd15KBed3A43nQ0@j:3MU_aTKUPZPeM?eB;FZhV_WjKFCO;jm
_X6gaZd@MP3LmLjomWd<^6N]FSA:J4bAi`i49_m=@KdlBjql6M@FXicjH=XZJ?A8
84\kR\W>`KVIK8bS;Lj_N@6lCDCbcIM^nK@l@Zab[UN57j[kZ=34GXO^@CJdI_>S
]CA5>:fYbk:EIa3:FIn3<jP6hQ7HQ05AK\S3B9oh]@cHYeR@4TiDUXheMmk7Q_KS
]Nm_Peh9[cQBRNNJL9kR[bL^P8lbcIM^c]QH>9Ph]@cHa^S9[:ZnBiMjH=XZJ?A8
84\kR\W>`KVIK8bS;Lj_N@6lN\lQ1O8_>DbCRINlaqOBo`OEllU[dPEm[GL`FJ5]
aZD5dIfa[9J>E=;n_H4FQc?hOJRmPaVC_RNIUcSf3iQ:kCGoLNDGZLC[9_:XnSF`
:]ZnSi5eV3h?RScK7L5i7ac2cRABF<1gIS5f=f`YH<Q:`knVO[\;cM1[9k:X\=N@
A]E>k_Gc:fBmk1]f9@`I_V?hOJRmHJOYOR5f=fTjNQSeMfPfl8U[dPEm[GL`FJ5]
aZD5dIfa[9J>E=;n_H4\Z:CNkJ=X:6W4GBYBq0R2_YThR01EcfChN]LT?3TFEhkZ
YPCoR5nq6McC708XdE74M?SJ`_k]BEVH<EanM@]LImQMfR0jHJeQ;fgbLKJRKW]J
7RZH\Q425=eF::9eN\a>^d=MMfTfE[D>4Q\JknYO0`FnIjJ1]P?9kTClCkW13hgi
>]Vnm;Ymo^L:8K?@jE74M?SJ`_k]BEVH<EanM@]LImQMfR0jHJeQ;fgbLK7S9`KU
4@enN`hh4AKZ@>3lbi:TQADE0j[<iAnq5<TD;f_U<G541BNOJmAdBcQD@A]Z7fZU
OP[F4KKjSRgcUNKQBNK5m4nT<G1P\XT[InN@_3ME?aCLSKF<ScV_4Oj6E5_O>kn0
6:E1KWL]Dg?WnnkLj1hmiLTo7>CnDnca@<FjbF^H4G551BNOJmAdBcQD@A]Z7fZU
OP[F4KKjSRgcUNKQBNK5:CDFG4>>MUO>T1:f3PDk4fdgk]oOGT`X=]=qE=5DcFKb
^o3UYdNmNhXA\=dFY\TWALOhZhBfTUJ;_];Y8a>nUK1giXoI0GCEVZNLD0hYB<OK
o`Y:P>IU6CC_Z0?eP8a[9oKK7ln8<fEjoij_n4oQU\<d3UN30Gb[W@a\E:`PMUIL
mo3fYdNmNhXA\=dFY\TWALOhZhBfTUJ;_];Y8a>nUK1giiXA3jcY\?OK]20il1`l
PXhEb7>Li9KJ@aJpC5G0Rnbca9[7]22TQ[3_0NPBeC8kgCb\7R38Kg]ge=l_hNj0
KS448bLMSOA5ORmh<1Qgk7A[LaiXhZiFFbhPJZen^PH7IU>2919Nld?M>KRAQPDO
L\aL?6QASOB5`9:ckknlVobca9[7]22TQ[3_0NPBeC8kgCb\7R38Kg]ge=l_hNj0
KS448b5c7Kc0S>abkknlVongOhZVCgC4>mG;9Klp6KC;J6E;n_5KJ[SR0eZL@18P
LOP2oBU0BbXXWPA=i?U?mJ@683R^a]XX99bfoWPMXDBAFE9\qAJMFj;FgZ6T8ABF
]GXg1]khR>[M2bICgceX:j@n@k7nKaj@d1ZkM61aS=03RC]a0ZjjFTOE_<oT[li1
W_m7l<FNal7FjX`Z[ccgZO^Eg9?lLH\?CeOio0ia=M5YG]_JbU430Q7F]Z6T8ABF
]GXg1]khR>[M2bICgceX:j@n@k7nKaj@d1ZkM61?KM5YG]_JbU430Q7ef>ZbFb20
8`AA8;]hqfB?oBSUnDIf7hKc24AP;1dU_`DFL:7;QZiI1dYa16V@QlnDTd2JH0`B
<_Pa\JnW;fnho>W2G\igo25cV4AP;1dU_`DFL:7;QZiI1dYa16V@QlnDTd2JH0`B
<2?DegCd_^l<ZVZUgDIf7hKc24AP;1dU_`DFL:7;QZiI1b<m4i<U@@b6jhDMgq^S
Y1f2i>b^RHEH:6m[mk^b2\G]F6gkY:_V;Vnm6hf`cjLlCcKSCX2GM_o;L[WiT8R8
L@B[i6b^RHEH:6m[mk^b2\G]F6gkY:_V;Vnm6hf`cjLlCcKSCX2GM_oHlG[i^MR8
L@B[i6b^RHEH:6m[mk^b2\G]F6gkY:_V;Vi228CV^D2Co;Ca92qf7Re>f>Ld8UF]
TMKK6eG4SCFkf_;aJO6X[QFDKmD64iSW\]A_S\\GEPHi12^ol_ImbJN:f>Id8UF]
TMKK6eG4SCFkf_;aJO6X[QFDKmD64iSW\]A_S\\GEPHi12^ol_ImbJN:f>Id8UF]
TMKK6eG4SCFkf_;aJO6X[SFe9<A]9T_^^U1Campb:I[EkHiX<C?OCl>RCn102mX3
IMaAmKW^^O6CYnKa4YPL^k;JC1VH0H>4YmW4TDSKG8c:nHdX<C?OCl>RCn102mX3
IMaAmKW^SI4U4l[``ABE]:E?YqOEbY>U\JgmPXHKQR^Uc_hhE9F1n15f12^l3@bd
jalOeDIb2hn^Sa0lNVASGYR=>BO9^Ci=\5gmPXHKQR^Uc_hhE9F1n15f12i:3I_R
8f:HA9:DGf=2pB`::fe2I9=R[^SjK3iDih;bYYm??@kECE:i5fB6;l^eInS6Fj9K
VpRQh3<Y@S=2`XFkdl0Ao]H2B2MA7V_dS8kYKYTYI4U716C:8UP@GcS^n7D;OS0L
OG@I0`B45c=2`XFkdl0Ao]H2B2MA7V_dS83BoN:5XFD:JKckiZF:pb:N=e?@f^`Z
k0@fQOh1DYf\JnS\QmKOeL5@TY39nTi_:80kYHRdk\`QQ9PbaSG0oKJHNh_@\UQh
6K4oF8TH5mZdQnHJWdCO]L5@TY39nTi_:80kYHc4PHWeafPI6hlEOH=eEJ@Lqc<B
g2l1b24I2[A:2=Ej8_F1k6X_N@^12?@ld5MdV\f4[_T?Wmkc5kkLS4cGF3@U=KP4
QhFN8LIndR^><;Ej=_F1k6X_N@^12?@ld5MdV\foJ4O>aAUTH:^jS:Ga3pei<d9C
ife`MN@JI:6EeKI0OkSmHD7^fnND0UJ_fPYQc`XMmgVO\5LSn@Y]MDNDMODS:ohg
3c5;NYH497=9:0IgOIHJTP7DN4D]B^o_fiYQc`XMmgVO\5LSn@Y]MDNDG7XSo]3g
lA]QSH?X:3qFZZ\:A5PCjo?8Z_7VaU_^LMD`Z`7C93Y^ZcDhYeJ7T<odX::HEQoR
F8i8:eeJJ6H1YQCAa>QCjo?8Z_7VaU_^LMD`Z`7C93Y^dLkU;gK\hGW]jAJnTHqk
=Tl1nOL\6a>Oo2pTUN<IJ`Y$
`endprotected
endmodule

