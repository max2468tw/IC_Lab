`define CYCLE_TIME 5
`ifdef RTL
	`timescale 1ns/10ps
	`include "MS.v"  
	`define DELAY CYCLE_TIME
`endif
`ifdef GATE
	`timescale 1ns/1ps
	`include "MS_SYN.v"
	`define DELAY CYCLE_TIME
`endif

module PATTERN(
	rst_n,
	clk, 
	in_valid,
	maze,
	player_x,
	player_y,
	prize_x_1,
	prize_y_1,
	prize_x_2,
	prize_y_2,
	prize_x_3,
	prize_y_3,
	out_valid,
	out_x, 
	out_y
);

`protected
G6B69SQV5DT^<BO`Z2n?4^`JjA<;fVje3F0AKPqCGG>_F]3cmUUh19<3fn22\2dn
QJaBm;bcQC`fAh>A^^o^\jD4lFpUQa<jYWlD6dJT2EK]9]GbeBd?P^DT8hlF[3=S
ZijS2N6RE>UMX:gTVSZOE\l?CfjoZ9<LW\qIZ6S``p_`WIb:XJ2hNaJdT4W_=UeD
<9>0EJQa]OB?4[bF1[q2Xhl^D3U9e1b=`=4;^HDfcGq07LckSqPZ;aoQMQ1[gh22
hc6_fCeb6O<0SlilMSW3hAO::91^]4p=1;852;`?YN9g;XkKMN=dT^UZgg;Oj@97
h96p[dCK9mpQFEQ2iU0GVi5BA<4f_<?ASTkSUeo2E4`<=3M19pKbWg;HiNDPQ]37
mh[GUJH6SbkF2P]3OELC\_i7qf`4ha=pPe[2=YAo53>U7U2bUcKQEZD1@mAA6o@Y
SCml[d9:T[ng<CqPJL1Hn06n3T3genQo@BdgR2@O4IQALm9j_Rh?g_nORNX56qcA
ITgF^GOM7E]Vi`n@Y6L7NMel;^_h6o4c^RqmnURH]8J@I6d9[jXb`T`m[W]UCn1J
88K2h3Oq@WYlUGOoHmi5IeVe[BMX<`D^k=I=3SiWe3lBHZjHWd_2KIqG4l>EC@1;
da>cD;dmck^[no`hRcc1Ql;1=iAqJUU4L83dO[0JQj06DLo:cU]>W@5beLWl7a56
qlQBfm9:o?24n`;`jNULE:Q<9a_2A2RN2SDf;q>4O\9fVZ^a@1>RAje>5LYL8ET]
5=76@YEY6a_dkBIGb<2I3\UJpV4UWUJ?bOXU9W6][K<Ia77_J7ZnHDc5WZiPRqX<
Fnkep^YYgN>b:H8CFlkdSm6iO549d;2C0m7bm2688@NJ:cGXHq0;^MDi583gJHPT
Q8Wijo=VBYKLAjKTYD\9e?9YIc2oGN@0?H0gXGFGk5\FMk@>Vq?SE4UEET?8m\J5
1[M112HX08nHCA0dV?daS;`MUgAShEpOfMYP[`17AF=ZDCPQ>jSjCDNShNIR;kFR
K6>WbOhCSj5pBfBB[:C3nbYZQC_8G0OJ<P?[g;Wb=kIlPOWVSL>i84=Fq<5B>K5a
bT`4H]6J8cN3B9<^n@[PTDmm<`TW8HSM0^8Rfq0KYa<Z`fm7^o7K2TK]?fnIkCO\
R]__`XT<FZWbE[`:UDpTi@9AI_0^V=80D:;BVkU51P>nTdoTO11Tdq8[Y7@D9`U9
1laXR_BcgVLQ8j1JFb`hMNZFgOqO?gbh<YLlEh^EQ@cI?ZR1eejNd=2pYjmM2@aH
?;a:M4Bk6i[YLULRYGY3Ea8lS>J062Cp6j[Z8NCW9ZCXS4GPkR7EUYW@qGd<ognq
=P[H\X]=@SCTUG`^TbU28F4KaknFFa<_l3d<YP6^cW5P9;^De^bWOieW]TgfGSf4
QWcN5aR7O5S15<cd60_B4C6ZnKpLRlb=EbhFTRe22m7GDk[G<_Qfd6H^BG6f9Y?A
@7no>B0<d^ZY<dTDQ86P[YW48U58BdndNmoe2qE^gjOh1Eaf7jB9fRH0THkXO_lk
9lU0\eQLTM]>P7alFJT2pn>bD8;CJMH71k?Am817QgDHh]TIj2M^^2OAfp?>hhMC
mB\\oB]nUn6^E3Dg;>daHo]j@P:`X25[30hn>AF<g2<VCMlA:@P1I<gG2Dq=V?2J
TqcggjgTqPOabEaW_=NQFQ@S4kmUDXj7NGGUko8l^c2JLTmT_bC:l`?Xp^bX2f=:
aJN4@6`NJjH3?1b:q>hKZkSp\j0`?0p]UWGX;W6U<W:m[\i_O6iQ^o=ooKW24G42
=_n:VgbPOEBIMDiY\>hR72]alqg@3c]0]DPg<d1YklbKUJdjSEKFbjfe5gM9ERZ2
1MESRLD3j@MSCU1JM2K6Y_hc:Ep`ba6S>UHR<GCW8[RLZ2hb<Zco=Kq0kUGM1G:K
FNQQ:5]c7qHcg_M7eBV3Eg`SV9PR[cncbQ8dgb_>5MZfO1Ae9[4SVCD:Rq8W;DfB
59g_^4laX`i]eMbdmA6BU`^<U=FLT36<o]nBf9?HgpJQ\9IVXnj9p>BSY_OA2F\[
ed^M6cXN]^nm^AFUSMcL>q\Gk]h<Ul6oDU7Q9;`aL7qhnDegh74LUA;>Zh<6IMT=
:gfZn>GF@D19mq1c9TOipUTQHP=K9]VM<d`NB4Y;bV]k^2<;CTL]]?2imP3jk`Cb
RV167_kOG;JM^<\8Rm0Hp=>=H`5Xc8`>UQL_Ke;e5_G4ml5[nEJg_5b1Q3D0KAS<
oNH`2kFWHP8Nd[]GkWF@i=YQ6jQoQ:GgYCll7lQLcg]dU:PEpBP20D0kK2lJCdD_
2>KLoeXM;SjcZ<;Qji5j8RHb>SRJ_p]IeAIj:dSWLaiY<`f2LFQ<O?dO]VRZHDCT
X538B?O3nV=fHX?=43KE>4D5qg@d[aSV;\lm9<]`f]`7WVXi;ean_`=ojQ2F>EjF
5gnojHM]hOWoeO_Gm`X_pZ0\R:a;ggECLC1aqTCf_1=0YndiX9:56?D4?o]DnVKk
kJO=moWI;VBBC:WgnA31h_<kGe3>1fXHUfa8Rd_>Wp]I2Efi=V9\m6KUhcALli]6
bM@R;JkXZILo82cgPD3aeXHod9Vdi]GP2^X>\]U3SXj5hUpQ`^36IQ\SWoXPj9L?
U\g5@[CcYFJ=W13U2aFUWXGnlI`6fUoY0VV::;XDGXgZ7e2mS?UqSD2In\SblX9E
iYmiEah2kXWq[QC^Z87J_TA8i8EXO@??ddqBhTN]Jh\a2f`dl]pUQk@_1`ep0KPe
7XpoT_6Dhq=[Q`9EAH5QVG@2B?=m9CcOYM5glXJC2HpTb;E2aDqTAaEPM<KhLP3Y
6L2]^bUZM0GVdXCOWdH2apZH@BBj_XeZWf5cRgoSJhp]\ZoQc1qM>d4Q^aB:Qd3A
219:;KokSUG0j\TJN55V4X^J[`:LhY9pCY2\_[o[9m[Kh:5^?OUlKS:JDTUcpU_g
ilC?[NP\Pl?KO:MI>pnT:Ea64qkfW5dhp;]Fi0Vq[k^4gg0k2Sm0BV8`2Ih07?6c
8J<V1CJJa>WIGYpGg@;LYLne9aMelBQo@5dPhV49g=Oq9NWl4mHZ8MX?[hN^^=J8
bPeOFPkggEOcBMN5lB:k7C3?=I80;JVqI[8E[\AFba3YdjIK>lAh852cp5f7C8FH
0@U3_@P55XaHLOfFTmD7QKIplH3^^>B;=[?`A^:KnTGZJ94IHCUEFkF\L=DpIl]D
TUgqW_Y<g>K<d1<K`R8<0iYL7kHhp@>jbgDd?^:T>AG4_ZnX<YEZh>e6`9D?mM3d
pP^KFRC>96cJjPLkB;mbDjDdS`@0l3jEG2Q`DHj<0Md;F;6q9L<CSm2pWI\HL:m<
1]^PPI9[02cq8EE4X`VpVDbYf8VV^k>[;NiBhgMm81DF2TNXe:mF<i]oCbigKP_W
=BWY]AhC7iWnmOSKimQF8V\NaJOGC7fgNNOXF`A1O8qN=G@1E0QdSoA^4YT4=\Oh
0Cn1\>gB3La]BPd98k?5JCHgbj6\ae0i?KTH4\^cDL4^]1W67WVLEfbNFXNLJ3RR
02qW=9>^U>afFMnS=9=;mN_O;03U>j^3fLOO7jUOjWPZD_;:5eqZS?Tm^S6:UP<A
WE`4ODWDEQ3OmCT3TiU=bJ:C8;FG^fhB?gSmVkSa[oj37]ln6P=nnqI4=33n@7LU
5i9UTg^T[3Ioo\f^FfMRgo?gS>4h`LHic?1dSoR:M@]R[h@l;BYS3kV?8?LoDEZR
Q<=P4^KT8f:^7Nd\B2BUYHE9AoN^mMq[P_hSHfQ\k?Qh7V=T5kn[M`]fFV4I0>h?
INRJD:WQgo3jG:RmgVAU:Wgh\eE8GV=1IJI^PD2HLBf8m5oJURNND:q`09QZg7]W
]_kYB9CR>9fVf1T:2hMGlpha4GFlca1QT\>hRkH7pmg9>>U3`MJg<[bfKVEB@@kR
oG20l:Y:ab?UT9n\g[42m?Yq0nZd8OSCq\O62EYE=Hmhh2Zl^U<V>oA4`USkOl=<
3dj^Y5GXQ5cSDEiI=i[?F]80Wp_76_dAeICQB31hEU@QgIKJlW0Vnq9g2gCPSqUl
N?`K:Z69pmB;WSnq\SSEK\3Y8cLS@]cm^KjT9Ie4Ifkd`D`[a31aB<ifI21]iH;M
pZg@B?kpO[J29d2<CI8`@<ZL2lQ6\fj>b1IjSI>G4Up_0B`jC1I5KL66QoIY2<JP
fl4Ck11l8JEP7mGBlS;eGjGWPC@SDeXA8g9fBnDjU0]RHW:hAiCeL<G7;4d?7dW]
mapFE<Sj_9m>Z_LjaKc=V>6fU1gi1\Ogi?mVlTe4622N7F`\`W:6g41i2F5[BZ;?
7;XFci=m=D3n?K;L6MXgVJIoU_ZiM<<6JVj5eLQZNq9:4D4k?;Y4gPiJH6nJJbWb
2hMFIiESCga]ogkl`lL2cJLj9gSPW4`]d4T3FADfTTR8ClG>RY`4ZJnN5S_7M=K@
Cq7j8c;A5dJa7B2fe>MI78oD@30opd?FdlXKGE6pnAXf>Vqc=1ILmk_IE0@0LRkU
BaRf1ga2\Vq[Y]IU4F;BFCU>4fZJilE\g_Ji@9MO>q9Bhk^@qn^>YQV_fm7^_AK8
602UUD`?f7i]FDW=L_N31Pg\b8DL82PafMS<4]Jn_\H7m@9cc@]T0K8FCaZInBMf
jXj^R6Ie7aaA7KY6c\7?WH9K0:5aEYn8\O[_:BOWbD?F?HonHMCKPH1p]hUNk8S=
kUO<cf98`FclKK4BdG_J[\8b<Z0:m=AT?`oATOAYNVFSJhT?B1^e28=`fH5JOo6j
nSm=Nf[7P@o`l;nQpQEE:emq5CcFaiELY:7fa9^g68ff\7DYpIT3Q;CpG^Ln8GjT
lDI6fd5lf=C54R]5F1XjRYCE[^?BhGH@l_U^jkqWBJP8JY9c3i]o3[4;17b@HS[@
[n_E0VX4Y=M``H0`XL5hU=LD\A9NKic[dJRW6=o[k]C_Q?7YW=W@4V3S]hMYGIN2
2n<XaChpZU0HgJq]D[YYJpDFh?ki?mI8_dhhNHUaL5O[[JT?^b;UoThn4I\m1jQK
Nf[7ijXEjjRCkS0Vld^GWil0;dR5GLR^ST?ea;f`RX5<0@B>U9S_:5d]7YjLGQO^
DZPOQbA6gLH7amKMTg5K\I@F_4Ohq79FD\D^Zo5M<XJT>CS:NoX=43YU8S?@5EKY
o]0K@EORKVdojm1W;<L]LNG^hqcne<BZRUVAlnhfcaAUKF@n`k>iM@G5kInRPmW=
QKUaMgEOK2;]23<9le^i<jg8`a40eZAkCg=o`@?L_?=?SB]\jI1LL^MO8lfF^]<8
0OCGM4\n`_c\9]FdbGEbJ@nZ4kahJO^5_SjZ04R6l8ANbFP]m`1>G;T:Q>\AH?_8
0mU`N2qL<WH6Lb2=\bB8HmkZ==9fAh?`AE_G=@hA88VPVSG=<k[?SCVbJSO4;mbA
H[EMG[Ik<De;ma_R1`T6AElLVDMaCPAhSl8?WKQDdamINBW^m:J?SCVbJSO4;mbA
H_EMG[Ik<De;ma_R1JT6AElLVDMa9naATp2YH=9o1TjjN0>6n>2@LI@4N8R@^_W^
bq;4J2nUZbYQLd:i2@RiVNf:]>U@`3ZWA`Ri_maP0dLcqlQ8Ej3N3OR7Y09><W6<
Hq5mc^CHC5qM3nk<Y^HbiBZcB63cMnB0RH\DnkTA3]q6Jn4C8Ul5=n33CE=gn[MH
^Cp^nEcVckl??e<Ofj?P8PBpRmDoe>Up;W@m[\R<kIqk]m7]Cp6[8>=adoh[mJab
6kl4ZTh56PF9fYQ4KQfkbU7eX6;oidjU4mTAHhCnANqTa_h0kPWIS_7[Hm>qSohc
nHZXRIjd`h;PP:pIRU>680KZ>S`c2:J8F`KCJZ4W[p8[BV<F`T?8\4\Y?NJ1^UWN
b8K[O\C``STYU^2mIn7SfDna]4LnfXkT7N[@:mdGR:=oe=Mm0ZmEf`5jEh0OF5Mb
jF:4a7ko\\>aPX[nmb5i>jXDE9A\h4IYMeWf2fmF7cnPM3pRcal4CcWGn7VK]dbI
[DUccNW?lR2BV0lFf?dZOC9gM]jlaZB_O<b0DLJcGDqMM=8UEpXY?gV3PhIVET5c
[h>@j8FA2p\61\UEa\ROGg5[j2U3DX5O1<qFCXRG4N4i9S\]j8C5e]Hj1OU4O:?:
]jplR\beSWiBTilY>mSigelCBEGqZ5DkJJIC_Sg2BV7XcWB>p4?[_dmldfOb\ho]
S5J]<QXfK^=n^cS6QbcW8lQqSO:O5Dc2@e>2cCd1_V8E4iY7KX3Z1=RNj9Mp3;Ib
YkJ@MmPQ<OiO66:ifU@8kR24`nCd:8EVcA_DCnZ3`C^@?4bao6R:WLXdaUNWCjaE
g>\3O><L6ZfUDN:X=RD<LoeGK[3<2Zd^cKZD0i3qSLSJE8qPl:fSnq?EOUn?q54A
G9mq0a_4HPlUgk[QCFBlgC_U63RUolUSdEZlF[iRWHP2J6L4DGEB@_aeYW<SeffQ
UK^5_ObQ7TC5:M]@Nll6fQTp\Zc?8n^:09gKPTVFiLCJ5mM>Y?[LZCjBYI77439h
m6=PjQLRbWXH5HH=VWmJSeC<lLJD;1X1@;>Ma21_j]IQ]gGp<b9\8GXmNHhcMEfh
06P:@PWnXi31eC`oL1PW=EjnUb>6nn85ikbkNCkA<@>[OCB`GlqQakORc0XkUf]F
nQQWE71b5lgh_d93@L;9?eD<aYme4[m<m`FB6MHXClDTNkC^l_7R]pP3NZ<Xni@\
Yg0Blf7]cK@Xf:US39D]O4T8Che_QYLP4e46C:gRX7GU?J52mF421=jEfK?m9VLE
h6EnnbX;<Bo1GD;8YS0T8;6@C`Ob\i59mfV8n=4X6lbl375HZFT8d_J_k5a]9Pik
[Pg[iYf]O0o>fmV69qKamGeh^V8ZWS4GO8hO26Vb5lZ85Ka?0QARVGnokcfgahCi
\W=07Om]20B0]PCAE\fK3eXm9]L17AZ=OZ>7SFIIgpjUkbo3^0_@mXJPbG_]YcP3
k2ZSUiB^pFJ:N[56SHI56HQVpQe]MS=^V[d@Qe:2ooAih]M43DhUjf;A7;geKIXS
=3M<NSUjo]M4gUF1m^lq9<U7?3oQ90BP<6PJ9Y<epHnGV80XWp]lN_TYYE]fHIae
>7eg38q^gkEC=QZU<PUONTY9Ue5Z^?M194@XW;54Zb40CpH_<Re4\0pm<8R2WicH
C1\^oND?8D2ED>qC0eJhJB[TOgDDdMRZ4:IAgAP6@iknXpDPJhcB]eah?V]Dn:f8
9HO4I`^GgITAhIoUO_d]U4k]RGOD7qWDHX<302p5<iaSi?qk?VI`]OQX[018dl`n
A_KS<>AF[RC=^PF<e_3b\M7hABpQRE;aVW:DiP5oWMdh51I_]@5WT?Z^9WSIBbfE
hXbA`;oEPPed@hhoWaBRVhkAedKPd`AaZCeI?^n7PD23HhEMMYq1VaQJC5c`\`T`
7b9ZQ@7JPCH?SMhDM:2j\N85?F8f3U_Pm_GDgP4Y4OhnU8fY:a3@8qc;@`Fi`:m]
80jNZiaiohSFVPmFb:\MPjfePPlF0Fb904Lg9iNG\2]^FCdDO=Ae8ABJ?1RGd_IC
EJkmQK8e5jYoqN84;RUH]310E_DoPki6>UBBW^aiF2e013IaAVIo5k;HjA`5ZiiD
@GRY45fY64ddfD4X@b;hFCIV[>:Sh5hN:L6YpNmhUZH5NLdmB1KID:=[IQ36gK7G
NgOpij9?46bHHFk_=nPZUI8pdo@`P69Yq@0j5>bLmM^Um>Ea9jV4cXjPFfcF`ZHd
>hjoVhKbP<ZQZ4eFMWH>qTl:4a7M^qg5@^:AOp:N>B\73UH=pXPM=64pYgA2m8po
3gG>=qKIToof;a7VEFb376Qmlf6Ja\Ln9?kj92Z^@gSEhQ@;@4=UJ1KXaph[bGEV
d:OMYfIfHYmM1jV?K4L`;jSJpVFlE59TEhIJ\6m5RYH5@5[HTGOX[CgEdS;IooO4
;?S?^79FL0RghS1N_hN`94KH<LWa2FRTVhIJ\6m5RYH5@5[HTGOX[CgEdSSS;>T_
NCN9SB9FL0RghS1N_hN`94KH<LWa2FRTVhIJ\6m5RYH5@5[HTGOX[CgEdSSS;S8Z
X2Vjo;HQbZ>aIq2[ae_g>a:\b^TXcM=Cj8QdkghQ7[EQe?\nTZXQ=Cd9C^>?AHS?
QS]0ZERmAbc<GdoV]VHV>]:\b^TXcM=Cj8Qdkgh:aVSU1m\j6]B0MN^J]PXoUgDi
QS]0ZERmAbc<GdoV]VHV>]:\b^TXcM=Cj8Qdkgh:aVSU1m\j6]CCGl1Pikbo`1G`
gRpkRTWGlIUKUJFR4DnQof1Un=Qia:X]fA4L5Oe34:WkI]E7EV3JV=2E1CMbTdE`
EHS:4=>AcIaKUJFR4DnQof1UnaQNd^5RKP7[?Y>0d9@naaZRNih40U=`TCGbTdE`
EHS:4=>AcIaKUJFR4DnQof1UnaQNd^5RKP7[?Y>\FA;37\8obLHjkBjp@_7\IFGJ
=CEddPm3=On[UQJA:5Lh1O`A<1B2=dcGB@GUdA0Sm0HYST:0PQ4T>O4@[aD[cnGF
=CEddPm3=On`KKif\B5\];P0<1Pl>lKMK@3kR<PLU_OL6TK^PQ4T>O4@[aD[cnGF
=CEddPm3=On`KKif\B5\];P0<1Plm[3>:cUNg6o=kYF;qfVF;P;lAbo:98H;dGIb
OHj`81KS<8l2`8S4Ichj8]e=e_9I0JZ=:nLC;>IMlllm9KELje6lmbo:98H;d495
9j6VheJ8\4BKR^bm70EjCYL`BD_JHGA\a8F7S>IMlllm9KELje6lmbo:98H;d495
9j6VheJ8\4BKR^bm7Ndh:YaRKWolQU\<>qEh2[JKDB7E>NP]UhbNJGVf_B^9JYK?
0Uh3Q`@^SI\>`>km@mNOD=VlA8Q5S?lYAUMQ\?\j55dk^mYSM^`?o4m^6@bn]ml_
OHUDlnfZ0YI5Xa>B=B1oiXSknDQ5S?lYAUMQ\?]j5DFF[gP]UhnFk<MB6<bn]ml_
OHUDln>84FTn]E[gBJmOURp;ObkjQhlI?M`QeXg5]iRd\D?:_<3CAGUkPPXd;K^R
]MAgU@n?^F2A>@dIOkc;6XA;ekO_VU1]J1mhAk]5]iRd\D?:_<3`j7@DS@QYUGFH
SZ^KC[HC=TARYQ^l>\M6cn9\ekO_VU1]J1mhALniITo6d=?]W[<D_Clmi_G31g[0
Ee2il\h?4PYqdAKXe_O\VU3aVZhAGhf=VX0qdUGFB`EW:]8f8C2H]JQ`_<:[hjie
cDCo[n1CjcQ9bL6L;lRAWPH666HLY5b\K68ad\7<A;4bRDin9oTgB\Z\]M:[hjie
cDCo[n1Cj^H5lhW;mOYHN14CQ25aI4MV6689d\7<AV>eI6N>hHF_]JQ`_[>Soh_G
XWQCkA_M_P:RcfF5ZdgjE_B5q]Wf;cd6UJhWQbFJn2<hK^jNjS>hcShf27n;0Z?m
NhFP@4WW4;Cof\mT7h0Yl\1X\@fDFMO6CJhWQbZ_^e]G`A9ijYmo:6L;H@Y;dZ?m
NhFP@49H<5>4@42k<A>CQehoZ]4S;f_9Uh:P4DX092<hK^jNjH^oC\GmnoE:iaP8
inU>AP8bBN7[DqG;GDDT6gin:J9F60]bOU]9:g?JX:G:U@]85Hn\1m^?aGd5cO?P
\0d=\N4[\cNa9AL;_ZK_6Uin:J9FHLf9Md\GIOR>_MOEi?XhMH6h27<PaWd5cO?Z
ATV=\NHa1EWWogG\;`fX7TKMRTH5J1]bOU]9:g?JPPOEi?XhMH;L64Li5LfNOXNj
b3p^BkV^bR?6Tomki;7MC1PVI[od3F2UCEM1VSfPD6WPbcGdC_8dSPlGY_k2Kl[Y
j`H8gI@?nR36Tomkif7OC7SG?SM2C2D[CENQNPoNh6N9iX6cCIY0LPD<gO]EA0BY
;0M^Qfh\f^_6Tm@F5<HMC1PVI[od3F2ACEfQNPo^iHRK42:_XQlDSbiqHb2H<eM`
:T6dNhL25MnfEgYZ_6l:1Ia0MO[]`VkOE@WBRJ[E6MfX8b7P:>d\iHHk6K<][3MP
jT6JNhL2B]PVPmT<RIb_4FK:>l?<eWjYP7jc44bZjZ;=8b7P:>d\Le=2H?8CET02
7G\i`W661Mn@EgYZ_6l:1MKB>l?<6n2[5ao=Yb>6m2lopf7DH@l82kPTk]I:54SS
PaHAA4=g\h9MicZH7`Yn<S>NoCEZ2S7XZ<5ol_PEfSXpA[D_kR1Ma[nkk9iPhX2<
VlYSmJ93U0P71I9?3Z:;2Jl7@j>]SXoG7H=6?O\`[Q9YUTa5o71Ya[nkk9iPhe=T
hj\Y[]`hcUFGi[RV7?gB]cK<a9=gbZ6ONL=W?O\`[a`8AY\S=CInbm4`Kc@joQ0O
VlYSmJ93UGO7i[RV_1baSm<4JenfJm4?qh6loXBdcJ84T;5<@Q5\Gg0\[DVc1?O9
i2oUmi:MNdO9=b:n``3jK?SHEfl1Yk72_lYO^3Kd>J84T;5<@Q5\GglI7_Vcl@=g
;SoUENJDgJlUi@On]`1^j:7Q=4`1<k6<1hB?[3K`Y2DeB=5j3B2D@BL\JDVc1?OX
im8UOj79j=M1SS04fb4T3qJn\K?Jm4^Y6U8Z]3F?Q<HCeWjZYNL3?P3M]5WF1>W>
I?l`UIfQVN?>SUZ9ilYWo:L?WUg<m[^Y6U8Z]3F?Q<HCkW7hhjo3?>\:bWmD1dW>
I?T\L[U6U<UEQ03fMBkOmaJmLO:@^jBDH^7Q>]RX^ESL=^\ZYGL315j@`b9TnJ40
dJCT0@NNdgqF1oXjY8<QnT:X7Xc^5BifbmJOgT9g45kNeIZ:4T<NfMK=8DQO@a:9
A9V9MXDe@<m7WdimT8]QnT:X71?^5BifbCYda3i^ZI1OTIXE4T7NfMK=H;nXGnMD
6CC9Ml7078GFWZ<gW[AL[mYS71>X;3cV]CfHgTmgZM1WeI<FW^XK]OQXMTOfO0Qq
R9WeMe_TN0oe=H=LD4[9hLWH;G\[\K_n`iiIBH5O\]bBL]9QL?JR:G:N[]82:U6H
U3fWSQ_8J0of=H=LD4[9hNa^?8A20fXD\KMKBH5O\]bBL]9QXP>Z@OEFXXhh766@
h^?o?d5NL?ZP_aC6X^BM8WWJ;G\[0fPj`inG9dCal9YS[MbXhVB1qD?HBoMB95];
:5<1SS>l;4F@I8dSUdU_HO6A]SDjDJUHe`@G22GF`G8\SEdAKA=OedKK`[\B65];
:5<1SS>l;EK@VD3S2Dm0fGSTTSDjDJUHe`@G22Gb0`=CaEdPlA=OedUQO=:5nc1O
kH<1Tl=dR9B@h8dAWDM_MO6T]g]PJOm=jHi2fQO[Mp`0DLXD=d_MXXiYWJLBfg\^
Y4`l3<TePJgAT2hk?<>9Z]FN=kom99PnDkCLm_okgm?YS:QJ=2_MXXiYWJLB6GjX
LjLl;75jDH<\B9@1?b>9Z]FN=kom99LXJ1dLm_okgm?YSAZ>SR>]m[@KXD@d<l\^
Y4]8dETePJgAT2dgk0\KNSk:R\X;RBqYb`Y``bAM;TZ?@J19ibinhbI3HAQj2JRY
WoZBYDU^SKPZk7VYTip7i9Je<\g2HDGfC@3Id^b9i>b<Aj_72W8GY5kQYMHb_iQ_
J=9[GQigV49e[T@F4jkM;BV_S^Y3XDjfC@3klT`JM62<Aij:6]3@41c<e;Q<_i]_
J=9[GQi`?KFe[T@F4jkM;BV4SLQb1dJaPNb`[^b9i<IOYj372W8GY5k`enBc5;<W
\REBeSkq::mFUbF_A^6RMS>hfn4bRBdQE:S2`]59Q@mW;ULoS[C1VJ`?P`;f07P_
ZO8GdYFGiG>CbPV:1N?oCMd;]k3lKVYOE:S2YA7jkX6WGRZ>4R5=]J`PPDa9?7P;
ZO8GdYFGCXFoh6P91N?oCMo;fn4bnFY2E:S2`]59Q@mW0d;_h\0f:NRPa^k2qK>W
j7iZRofCj^eHY=]0G6BDLUjj\?<AGY`CbI;C43dDL6G5f>Af=O`X0XC8BR7Ki^j<
FmPAg^H2GemHT=]0G6emEUjj\?@\SkX3hcQQWG@]:^8mm0PUd;`XRXC8BR7KiE46
b<=AS^H2Ge<CAd?RD7BDDUjj\?<AGY`CbE>FdGVATU3O40>C1q[KZJYW`7IOB;]O
@ORT\nESG<^2:e5glj7j[c_if1@OBiFmVC1nLV3^PdnZBRQ2Ke=CmKm@KPP`4DfY
@RRT\nJ^?XM2:e5gkZ<`\^Z[84>G;=A9hCMkTL3^PdnZBRQ2Ke=hJKZE`NQ`4_fY
=XQ^DYESG<M2:e5glj7j[ceAT<DkOd>>j\27>OqaODe^<d399Hac:Y3_UG?g=2;G
]DnUa_Vdg3I_=eCWa05Y[[ZXh:8nHe0fRd`1DSeHj1aH@m_T3k3^:Yn_UmEg=2;_
]D6Ua_VdglS2LdEYLKbNGR1Xh:8nHe0fRd`1DSeHj1a9edY9Ckn^:b2n@Gag=2;_
]D6Ua_Vdg3IHJmLd0eE]o9R2TTCp00nLS2@g[=HYm0LmBX9CgbGB4V6E39<E8?gQ
_7F;ZG7ThP_mN9j18O\AV[LOH[SK8J95]2W_XcR]m02GNX9JgbGB4V6E39<E8?gQ
_7F;ZG7ThP_mN9j18O\AV[LOH[SK8J95]n@g[f\Bm0dmaX9>gbGB4V6E39<E8?gQ
jBPf@gnLH6c;@FfXpfHg0<gSg2fO19FSP[<DVm2d3SBRZmPEAKk?B6cO@]`bLh<E
Bk3X7q]<Q5bI2:U5kLUmC9PDeY6WJnBcDE`D@glGKhl>lVT7W@MdViWHgfgk4_8:
4BlJ98E;@0hdA_S;k<FQlZ=ZeJbWJ0a?DnjLQ3CMCL3O8YmlCN>[>C]3S[lX63]O
d78Xl5jFPMLn2QU55RFQlZ=ZeJbWJ0a?DnjLQ3CMCL3O8YmliGZ<m:1hgIfX6b]O
d78Xl5jFPMLnBQME[]8?dEKWaJWePq4>WJRRX61H0>1BUanLUXJRm6D]id;agCYk
]VjkXcFN:eZ\imk5GRk1aInPP7E@3QaN]@c;loih@mdC7YJLU7JDeMgPU_\ReGGT
ckGeCgSe1C@NbhKGk4N1WY95`7>5d3doJUEKX61H0QRaIOJLU7JDeMgPU_\ReGG:
8cQ:CASYWk[h2_fHb4<1W`95`7>5d3doJUEKJPRF6\mL@od7BB0@Qpge1b9dIQ_@
[f7jEd2E:OWFkULAmej2D:FhUIGA5=IJCEJ;nRgiYG6:h9:iiI0=9FE7=cPnFmY]
Iia`bH2EHlmShGE=BY>cMP0fS:k3I_I[7aYUa9NMM^=:CGEGk[RlWN:FT`moIa_A
LO4eMHWa:^Y?h]E=BY>cMP03nH_2dPj0oMBeWI5`:fLSajEGk[RlWN:FT`moig3n
7`n?[4BKNNPcRpKD1J:6Am@?QYA]ne2CJOZCE`fnBS<AlCZ9dR=fjAnY>^=]\XEV
81gR^6GBb<02hFE4B@cGP:\\IaPWHZHfR:1OG0g;1j9Af__O9j@ML1>hdG@m264_
MIJDdQG`m67S9i3L2iOXAdEX81bW6C>A[?WgE7>nYECT1c`O]VifjanY>^=Ykci5
<<9_LJdID\L?b0E4B@cGP:\hI]PWHZHNmU1OG0g;1j9Af__J69@ML19Fl2SVDgT@
<JZidRG`Q6>iK9;G\kH78^aGlpY?:[m\bCnZ\Z3oA069hKGKfl9XM3^SPKTlWli3
?QoTYZ?OH1F3hMcPpfaDF<3[RdI5IjN?o:1l`oXH4PjjWNe046XD5Q:<<@8R<JmO
8BSEVUTSY3IaT@IiMiC0`887BW9^JL5j3o>Q2Q:Y7ficTU\mAR_2@G14N97aV`nZ
=Q;OD:TEFI8YLnan6ZYoSJVV16n6Q5@?1\Q_0jXfnlWH[X_e`DG8oQ:<<@8R<J3J
Q<6J3Nlni[Xn<^gdSl[?\Jg[2df?M4C0T4j@<Nbcj0icMU\mARRU@jUnEAN::FB^
]AYKXGBR^Y=q\jEaV<\I<Td97?133MNA=6\X7<C_642\dU2DCP3?V[WaQ72WZ<Kb
8Y67`\fT0eFeood5^QUHaggm]Y?e2RV6_^DW7U7FCmG@k5XKhn^gOe1LH6M=N3[>
Q38<f:F2RN@]kG5ZKh<nOggm24`L9eQF0H6FIkV9<b83\15fCP3?V[WaQ72WZ\61
g3hk15Q[e1D<PlE6n;\n<LVDU>HFVYVHm\TFTU7WCmG@k4W8FkajjbC2hnkI`]2J
k7UDQYp`dL?AiE^\QgZiU_kThA\RGf]>IJN4<h<CBEjiCbP7_[cQkh9o\fFT3\OX
=P@Wi@Pd]JWcChaADf[k30kPmHGSO[fWE=e>YhmS=8>QSWjB>7NkXBFJo9;Ld7UE
1X@[W7=AhYmIK9:n\Md6eJUmmZ7_6:GTOQoiXE\L=P]iCbP7_[cQkh9o\fFSnYG5
5[OE2CCOOG\l1E;\J1l162hTCWBj0hADE=f>YhmSeWWm]eP@27<R2i2Tb>7a<Vh<
XqFdoQVP?BY;7CV^9gV603Ze=UB]?]l>SXflQMkZGYflDRf73YZeQV6SfRe[FIC[
TbXhY=eNTOA]mQlkoMjM_kfimH9>6]Vna9l032A:[8OGgWAQdnaoGJiP@K\Of3K=
KbHg9G?\0\`1UgbjihBZUGNU]T1Vka`[6gAbh_ZZG5flDRf73YZeQV6EM_\`KXTC
`dc5Y=BEloYQ=F^kOdV6aZ7B]V?>6]Vna9l^G^_Yn^nB?oVQDjaYQ7M;K2SkpR0:
6mk5BKJ;B[;Y8NGf_i\6gV\i:dNbj<<76734ZOf40\<k[8^\InNSf4eA;iOde?:L
5A>H4iYGKb2E^]Gf=kS4koYYlCIAi@`iNgG1i3Z>8GYAL`8a5MT\oj]i;NhFGUDX
2`S^dmG6>b;niQlXJP4OhQhldm[BXXHW=XjF9Of40\<k[8^\InhKk8j?>RKiKn6<
U`=nElfXMQPRPNC8E9eIWoYYlCIAi@`0_EFS2_hWi:Qa8]JYK5BNG=mp1NU9MAQj
O_AEoDSGSklO6G]6>Q<W^7KDE8GKd5Ej03Hp`0JjONZ??DlY9]Y@2dl?HG4mXDYD
5ml\mXVD7WcL2DhJ:Eo?6W>eT0nD=>:K6LR^O[_;dH3mBhmgK:6hEdlhHGdN=F05
<i2eMbgGE=C7OQ>4PoQk`W2h564hE51e`4`UT]Fjn9LI;^CKc=eD4E^>VPYmFBc_
iES7\15O<\PcPDhe:Eo?6W>eTZE7E1=fK2a1od`e2@F3hQdIm_6j26o_1U7E=F05
<i2eMbgGEa^BbVJ7LojE`8>^n]fnPmq<mB?7h521l]RAENMg\o4f7EBO^W5Bl>7Q
fTaIn=_3CHdGf;XiG;XATUm<`anFb_F;Q66ib?PO8:ElMQEb\oOf7EBBP]<4nFk_
MBGKbn@iK?X]h3>@GBC99T^T=B2D1og[e;RN2HoQ@h6^0dLYFc\838cC13JPbB^K
hCl4ho2i4:en6;;iG;XA3?^_4>7=kmb@f6SOkPe1lYR@MQ^bj=5dGkZBP]<4nFk_
MBGKbn@cieJ>H\hn]iW^=0JA7p8[]iU8j1A>e9ETo>\9ZI8\0alKY?SnDh7gG\9b
8H1W>j_alb^mKW;leoWib[M=N`]V_:hA5TcdX>YTo6\RAYINa]dS27^nM:mbdOSS
>Fb]Ya1\OWaUD[LXHHcZQia>NOYLBTJMa90DEUaCn@2e34mSkS=jZ0nh:LQ4NO9b
8H1W>j_D<]kDLGClejWib[3G8<lR408YiTfXX:QkGUS<<YchjpS[2]P`W96;O84G
4;O<_alAKMY_F`l[gm@0Q8G]HlWlO;8iKS38IL4XYd2jZ9?TKCSFHmC54R:@3d?]
I]f=i@X7\e8X>Z]PgL:Tcm94`_I2mR@X3;<He1R<Xf23DhI6kh^P@3hicSPN32?G
5kE@^Ik2F5A]k:4c:^k4O;G]HlWlO;8R5<\Fe043Y?bBe9hCU7hoZX4:\487K:nF
kFSUYQXS6p32l3H2dcVj[C:KT@51mJ2@S=9\E;?eDIKUJ>=_O8TK@GiCa9SM`aXn
2hkcGimB^5^WA:Cid2Vj[C:\5h`c521ASZTF9VSe42KWdTm?3G`Lk;3f_:TkF7?P
j7UkQEf`M8DWU7n\HanZ?NehG[3jaGJCbBKcCCQA6U\WJl=_O8TKSKGFJgSX>RnU
Rob<`B^EEP3WA8CiNF[]eac?bbEk@BPSDp`[Q<23ZeOBUemVQ9f3Ujm0ORZB0o2K
o1hJTjEhmH4MC:Y@?PT\4<LlMT2FiGglKjj[R7ifZCOBUemVoDnLLG^POIZeDCg4
^jhJTjZ>nnZ@M]_ieH]cme[CQ04><WfCIi_QN5M`TL^UE7o?6__@^KX^U`66;fcT
T@hJTjE`@hOBB8k@?ZT5I:SG?52:OlglKjj[R7ifVkBT3YiF]SFXK<=_@pVkSU`U
QKcaLTOnGhTFZDMfcFi<4\;1V3CAR7^3lE1S:`^8<WB:oB:RmKdJENEWZBb>Q3[4
QDcaLTOnGh^MiQ`7Y=<bDVP7H6CAR7Bl^mCYh<ABkFY<:8]j^@hENcR@?L;6ZQoF
oJc6<0bejVglobSW:\7?aUS1V?CAR7BlbhlIm2^8;jg:o^:RmKdJENEWZBb>Q3[4
[S_n=g\\:D6gJnO9:p7C@jLfM_B5Rg;P5?1PVEecK`46CF<PQDbCFLTKm^=Yj1O4
5NaD][nG>WCEEiPmR5OnUWKiMHB5Rg;P5?1PEYcAKA@G]OSCQd_O\^TK>DQ4j:O4
5NaD][nG>WCEEiPmR5OnUWKiG:5L[eO35V1PeYlK0^@3dg<PQD_O\^_I9]D[n`kY
ZM>OJmqG7c^G2=oXbG7\DKl9ZG1^9hJ6`nCKCeJ`PU:ORYmi6IiB6[i<eS660O]5
<m=bd^77adCjJ=mX<n9KAlS@gaVgDhI6`keMC@I8]\jH5gii6IiB6[i<eS660O]5
<m=bd^77adCTP3nd9bJeDK]9ZG1a60bM;F6ZC@:8]\jR8LkZjJ8`[MJbiJLp_n3A
2K:oNYfTYa0S=Ap;O5PUPV`@534EV;5EWT\]\joAlB3VVj_66JTf6i7A3ncSCdbV
iAAj^5j3U[6T\A6a>E3dlg3oUJ\d=^4S1RJAX4YeiMVjQnBXlHG1DC42Q?R0a]VW
<T_EP448d8hib^ja>E3h3V2@534EV;5EWT\]\:[6MOh`=FAM<nniiL1SU\N_CdlV
iAAj^5j3U[6T\A6a>E3h3F2A1fI3Km1j?2gjVMpd?Z1dXdkd8I3eIRRGPGh6JO9?
;1_h1\82;;6o<hO5S3A4D]9S6TlU_;e:=9A94NAfWkM>g>4C8TEg>2nTg@nNcY]X
IGC8?XWeHmJU\gd_JaO]0>HJh[H95e6MP]hdSjlfC;bXhdbd8I3eIRRGPGh6JO9?
;]JMYjL9HCUC2Fo@n3d4D]9S6TlU_;e:=9A94NAfC;bXhgbK;V<2@:Oj01N<GLp1
?CT_>cGA=GZ\AgFXK9j=VV20O:]LcVUDZ\S5YJBPgPeMO<DAL@RF\j]V?<[;`ke^
=767D<oK<3MNX<>^PX=aL?W0?ClLiPXPbM0I2<Q6Tc>?>jP3HPAo7HEk7PR]0FNZ
E7F=EcYA=GZ\AgFXK9j=VV20O:]Li^U@Z\j56A06gPcDj]8CC@@F\j]V?<[;`ke^
E7;=E3YiMTQ7g6iQAgG4BBpHBnM<VD5QKU@]f8ZZMfb[lCmKK:FgYnSKcklkVmYo
nOFWON\;1dmQfXl_oA^5XllN:J?]\6iN=nYRG]SYaDl[8TQ`:FkanUQ5c`lRjLJ5
g9kH?P>U38>Ta<4C4g\S_\`7L25AEDTQKU@]f8ZZMfb[lCmKKFc@lPGojl`kVmYE
^P?>KJFOehJ:KgZ_oA^5XllNL2_AELT=^`nPM;Io6]6WXhqV@I4O6LA>hC1OfLX4
QS]nc;3d?QXjcTpmN@LoG_HJ[c;ikHS6^YbB696amZIbh^c3mTajLDQ3n?DADQa1
[<U37M<PRIRGKnk>MPQLWN32IkfKQjCA4W?;JBEW>2jbh^c3mTagg_60nH@4j[Eg
2QUiN8_=R;G30n@Pi>==^XKm@BW53M]AiWZ4VXm7TODQ6NZd_RC`^P\1H^_;`jlT
4>XBEhc7@LCUolRmTGWE@`Gj<cmikHS6^YbB696amZIbh^c3mTag^PG11ZG`:Tb_
UXj0CcXd`phD5jGYQXTm:F>KlP=:KRM8WI4M]``K^=hK2OoAI^EmkeO[i8iC<V61
gmU=k7i8WR8D4e]3=5eWJE8j=H?h8h:DjM6mV0ZG^dhK2OodK4Qhl1M;5U1U<g64
[5Cm_>L?2Y8GUQ8oC1:PJ08>X=2T]QM8WI45KFWj8H9EQfa21H4>n[XGD`fCjQha
B7`mT@i4K[hnGY;DLZ[`MaNa1f]9e^7l0X6mV0dDbYHScg?OQbQhn15eG4GX4]LL
2507SZX@Km50VT9JQ8Tm:Feg7Z<6PW6U@>^l^EqY:LPNJ_T[bS16b[Jd:4d@ECc0
lPJVQKC=M4jc3iTJfF>cJXQg`fhE4QXV@cn<_Wh:8oeDH^i45Zm`Z;DASYIA\bM=
gBJF=KU=M4jc_m[>?9k^]f226[iB`^jQ@>UW1DdOOn:]mFP\Md0CN0^eS@S@ECc0
lj2c\<[ckM49bTN=@=MCcK1gGfoE4QXV@cn<_Wh:;cccF4[`edJf;GA\T0Fk6Vjn
j284K5n;TIMdGPO>?<]j^inD8AlbA=4cC5\hGJ=6RLV^H_S[bS1RARRK9\[R1h=R
Y6fqN?hPVI]S4XSfdXITI7_2W0:6@[f\_CEXXFgUfC_g3XTHlXLY38IANTZ_]\J4
9P]?oN2f?hMB^NcVUPSTXHbcOCA=3hcT?N?g_[l9EkES18\H[6LLhkj0YAe;mGiO
O;?i:\JXdk5HU@06I??3SkbF<0::@[h6fHiP[MCDN5m[\V<G6jAe6011S>4I0G8c
MPNPBab2`H;UXk5?n@_M\O>cW0::@[f\@NF\<POh0iEP1gQQ;3TXA``P5C>5jIUh
mN;B\VAfM4]S4XSfZlHA2W3:8=0;ebU2p56On@@[777?:T]c0Za9T1bZQ3KB5RAZ
:V]C8aUT3Zo39ObmQ87SQk@f[N5]CWnV<_K>D2Xj82AbAkeNRnH\OT[OR]b:D2?O
C1[aXoAYG9EO7JK16Gb_Ok]fIU15Q1IeZ?Vfj\B488]\FGdYGLQ[FM2O?]`j=Nf@
0>2?3C1TNZo793F95Gb^OCh]HAO]ZnI\:K:nH?Xk?W8?3:e<;naj`NSXDV7H?2?O
C1[aXoAYG6=Cjebm@8KcRRoQ121jln[]W8cUCGi[\77?:T]c0Za9T1bZQ3KB5RPi
K_bf1XBTT^@oFICpVVJn;<CP187_?lW[C`G\TG<anTUYgof;S:UZo;O_CNFi:RPG
lN8n<U16HMFi9GN2VjHL@AF;cNP_BE^SKEL8CGQ[2`9T0IlEAKX]6YV:eeW[h=cQ
0Njneo?ClSRO4Rh0F]in6b[SYJ0n;0J>bnXH2875ZD4f9UL:gWH`Xhg?6l02>1Ym
An6a92E\?PXmkT3RVjHLMWFD187_?lW[C`G\TG<anTUYgof;S:UZo;O_CN@i_;fN
VSI8LKSoKI>p>C@7P`5EkeXKYXb4>4H3=kOibdA;4>Ck]>RFj=aGR2SnAAbinVLG
BD;8c_bBaM]dk8BdT<E6@OFKf]5=hgH1Q;J;e_nl;a21MC_2YJ8Q?eLgM]P0j`?I
mQYARKANJ9hRHZAjO:LB1lF3\iJa<lElgR`JUUZW:U;_d]9m18:Gee3:hdgnnVGG
OjMSLeeJ89DIlL5@ZZ5akeXKYXb4>4H3=kOibdA;4>Ck]>RFj=aGR8jj2j?HgY@b
0ZZBQDqS[28Eon09YfUE=ZMN7]k5an3jno;CF\NAlUZY5J@Y^Q?aL8OMaNoWC=f6
IB@JUBWb:FiMIaC3;A1NBCbJ2Hm2T76kHhNm_]d2;bbba20<bj=4Zb`P^@C`b=5F
i[[X:UcXG798CcYi?95NFQEZdaJQ9Cbb0EkhfdYTO[=D>K;@o>JdBARMaNo<Ok>J
WgO=@0UI\mQQ=nj9YfUE=ZMN7]k5an3jno;CF\NAlUZY5J@YDg_0GbD[A66THno5
Wp`<UoO35kR?2XJ^ZZU[9F<ZQHNXjjh0Daoc[d1]6``bUVA2i\WVHCDa3f9K8V>6
Ralkjheh@f919Nljl22EXSPN@PKYgh=5MMKPLNBP]ZBXlH^C23\<AiR4B@@n?Q8Q
BIRL[9W0C6P0nY>j8X\96ACTCAbgIJY;75e8NLM1DfD4=h2dSkRVHSD7FXbalRno
cA:>\^bP5WR?2XJ^ZZU[9F<ZQHNXjjh0Daoc[d1]6``JRaGHG>a_P4KReDG6p6iX
jLgP`kO;;X[QRJm9gnBAM`3Y<qJdaIK:GV=\oOe4oc\?m=bS@NM>A2];`c>]4Jan
YFX`oJbMfMYHB1ghCdA@Z7BnP]jUjjBKD;VIGgHEKi83Wm]HA70j@Rb91WC0m6CA
3:WPe]d6PH]b^JYYjSGF=Sc>N`CUU2UaNoT79RjEKB8FQ1QbJY[:E2NbYIADSW3c
eNfDHK^[\lV]\_Y?j7GF=S?MRG:SmDd;GL=\oOe4oc\?m=bS@NM>A2];`c>]4Jan
YFX]6Wh^2VfF@k^[E0ebq@@Z=>[39@\ZZWe3HXEi`llQANVEBMjGENlPV>`XX2d=
gRUO]H0\IK?n>m]?4W`EOJ8WESZS2\N;J?R=m][nHeo`\n6=gF[j6H350KjVF38J
4DO:kX_6AK53^RjXn=EN^m=LX1ZA23Re\XR=m]U5F@[=E=;7lEjbjk?jmUESZ3a=
<RUO]H^WQo53aRjXnl=;hH[i<o938@\ZZWe3HXEi`llQANVEBMjGENlPV>`XX2E?
j:o_c]6jUl6^fClq=j3IbR6`F7DE>Age8NaDEeP6L^SAXUN10LEm105\0PCO`[[7
J8057IVWWfU<g^3Z_XgF5mCl:PmA?SR7O?HCB;TR9KED1[B7mX5=EoXa[GFn>f_0
N@n26DCIcHlOS25U?F^D;CC5@11=QfR\O?FC4V7P_LidA1X[SROiL:1Q<_Y[`[[7
J6@9?2C[cHlOS=MEXU6M@E6DF7DE>Age8NaDEeP6L^SAXUN10LEm105\0fj8m;?O
<AkD18T9n^pRHd=41nSiNUX4hJa`2InjcmM:AQgPHD2[khfeL=j@L9;XD^L:Dl]T
eEE=_^BVd?292U^oL4:gGnh76m`18\0hMA1YQbnRnn[TbNbjm^3CHV4:^8:71`5N
69bFJdBc5TC92T=1cHlAo`oe6m21870YSg68NJ\`E6Me]lGkYA@kSiKXD^L:DAm1
k@CFJdB7Y_hTML;J8n;iNUX4hJa`2InjcmM:AQgPHD2[khfeL=j@QglJ0:]Z\g>M
Id=_=qBL1S;=D@]5Ik@mQMUL9;djEEdiNeA95>7PjiO8C9YFA\XFYm6F<HO?FGM=
X2BQfKEcB^fmHZZJ7]]:>?kP^R[Ej^^SHLgHMFU\`\5Y5FB6[?Of[6ZJ0@iHA7]C
VS\1UYPSaJ7jNSk5IQ@mQMUL9;djEEdiNeA95>7PjiO8C9YFA\XFYm6FYH^6aBS>
jo03>4VYF\:S<2lH`6E0hX?a7l4JnqDOF<[H9:TcfW@<\;0KRHF@O^IXX`?76NOU
31KSQHRJ0=Z=H<UD4cb2WTUV5\6>0diI8<YflX@i^\l7T3B@ai9cXAJNP2_1U;ih
>FcW?GP87a5NaC8N:F6HT_^k5kU8<I;VK\fBH];cf`@<\;0KRHF@O^IXX`?76NOU
31KSQHRJ0=Z=H<UD4cohNeL?LEORK>0`iIo5DE\no1B8hZiUXcBA9p;Xn\]dTPOJ
iMmc5FU]VY@RI9cIR7FWI]ASFIbQ4f9a0lJi^^=cTH1i`KkWFEGJ@XgmeZ[SLAY2
^9SF2R`BFUGeWJDH\mH291nW_]N1I=ANO^o3>^c:bMP4L7kWiELWW5;6SX@Z<nOJ
i=mc5FU]VY@RI9cIR7FWI]ASFIbQ4f9a0lJi^^=cTH1diG3a[Dh:4;3L7JQR81<`
El<]F=;1I[U=aqB3BVBbiB8ICU4cV<0nSa?K`QY_gmWij4cG4gI6N8939fd9^1Rk
N5aIL:^o9UT8LkZa`D3mpdQJJ3HCnKGV9Y;:EE8`3N<1n7o93jI?iJlKBFM=[jhT
2S2S`7B=A<=IgMEkEKVRc8]Z\1N7e@<`XM30lC]@mmNm<JN8AOL22cPjQZ]Po0Lk
KS2be<dSnO=XPME5EiP;=Ed3:Z`CfKGV9Y;:EE8`3N<1n7o93jI?iJlKBFM=[jhT
2S2S`7B=A<=nTdbbCN2^8Ed3:Z`KKelZ@N\8XJ9iGY@op^M^K6^P?]a>2\W7;H^h
YH0;;@mGja\e8O1YD[P2PL:AX?Ka1LYjMYjAm:5SgI3>D;_joTb7OZmX]7\7[fBR
Dd=_d^HZ[_1SWG_GHXa66XhaBJURCk:2cHWAbSHGdUDVM=5>c^VPl]a>2\W7;H^h
YH0;;@mGja\e8O1YD[P2PL:AX?Ka1LYjMYjbgSHGdUDVM=5>c^V`lN6]Y\Rl8Kd0
A202p3V32]k_DC=UCKRC2mKTA9>[`Kine75bJTnTZ:4MN0no0]4@aa<M3C<Ec]YH
EBNET347P_[9DX[W=7VC\mKTA9>[`Kine75bJTnTZ:4MN0no0]4@aa<M3C<EcCLB
JWHAAg0jClT_WC=UCKRC2mKTA9>[`Kine75bJTnTZh5WckBc<6P1eDL5Op>1\;G8
DaT@<JZidRG`m67S9i3L2iOXAd@PA:2J@I2NmU1OG0g;1j9Af__669XCKUZFl7SV
DgT@<JZidRG`m67S9i3L2iOXAd@PA:2J@I2NmU1OG0g;1j9Af__J]j=;_IZFl7SV
DgT@<JZidRG`m67S9i3L2iOXAd@PA:BnPk[E16F]aAd`5aq\PM9S]jY]5\fDgU`3
bjSiTD?C_R4R]Qf8HL36>b9cPHRl6]HcO0Gl]P<INEklHkPH5^A=\jS]5\fDgU`3
bjSiTD?C_R4R]Qf8HL36>b9cPHRl6]HcO0Gl]P<INEklHkPH5^A=\jS]5\fDgU`3
bjSiTD?C_R4R]Qf8HL3;ZOBKX57[Rj726>mpmZHOleFD4FKk2E6LZ^7Jo>nH[9;I
2jN0lFimaZdb1NVTeoj>XBF;5CeY<[fDde;bU9e_59FD4FKk2E6LZ^7Jo>nH[9;I
2jN0lFimaZdb1NVTeoj>XBF;5CeY<[fDde;bU9e_59FD4FKk2E6LZ^7Jo>nH[9;I
2jN0lFimR9R11^::mb^aIWOHT4q;kTCIIX@\KMKBH5O\]bBL]VknE8nOk:;[]82k
n\TR^?]?d5NL?ZP]iGf6R1mBohi0]KcOE05_KMTBH5O\]bBL]9QL?JR:G:N[]82k
n\TR^?]?d5NL?ZP_aC6X^BM8WWJ;G\[0fXD\KMK9d5dnoGU8hBLUXfj9Pp@N2T[9
0C>QF\jBZKDLT04=Ufic]<pf3DS3Z6[DQoC<DmVJ;929?@8Kk9=;Dg9gbna^h]kR
deB4HZO[1ZkLafhnb@H@N<lWGSVgd6[?Wh`8DX]h99o9?b8lGTB64gBgbna^h]kR
deBmnNeffi^?\E\n\kfXN_5f^2dLi6hDQoC@mm??3\Un^E<e@?<3YqTMTKQ<[?15
>TjQE]^Y9IGS_eRHVJ\]\]:L4:e4SfDiCVAjBWc]<CE_l;S]jFhnk9jofY^NFa1J
>RnQ_CV11DlS:Z]7T4\]\]:L4:e4Yf4Z>7FjB5c]<CE_l;?ojV^kVXTonf^WO=8;
1_kQfiKY9FGI^gRhc3dXE:EMU9fo`q9SC_E^5\K>dWhL`^?_FDQ:2d8\14];T\RX
OcCQbHAkd_AGO8OFM0ii5_Wi0[3WAS9baT>9BI:7c@D[?R?F9>FS0<8\6\UnGLZg
3A@^@Okdd_AGO8OFM0ii49Ai^iMS7E9ja\k^0JW7gPGE;0cfMfg:Rj8<>[lA^jeY
@Y<?_H>1@Uo99K2dqS<enJhR?fK:^X]d?dc=PUFe^d7a;R62:8n7MLGAM<4lD2Bi
l5X8QKD@Polie>ZR>^FJ;bDR\fK:^X]d?dc=PUFe^d7a;R62:8n7MLGAM<4lD2Bi
l5X8QKD@Polie>ZR>^FJ;bDR\fK:^X]d?dc=PUFe^d7a;R62:8n7MAQ38bI\cAmY
QTjVEjXp5L]3Y\h8>7Z>cVhM<]q[B<9Mh\6@6qVd=WKoqBTDDY<Bi@BP^BPUN]ip
3kfbF]Bqdk\BVOnZHc211\3PR>2ES?lmNiCWP`Q[;VpbN6i>4q0PJ]2IcN=TKae<
9G?bUgNY`d=XY:JoSRbC2TBRc87Va4e`;X2cl11b_Xd\S[RJZ_6K@6E^eHhG<onK
XZ2aGdGhh6YUM\]F2`bC2TBRc87Va4e`;X2cl11b_Xd\S[RJZ_6K@6E^ch=TKae<
9G?bUgNY`d=XY:JoSRbC2TBRc87Va4e`;X2cl11b_Xd\S[RJZ_6K@6E^ch=TKae<
cG=kQeGa1go]TJXiV4Dl0H3i1lHYp8Fk5Ii3Hk0[jWfRo`c8ldP@BJ[VAX[1?0[=
GIMCWUN`FeG20U<?nebB284ffjfWIN@S]]6g[bSBcdX?H3B7`WRC^S<L@mkh?f6N
nUam@I2n:TM4M2cCngGBi84DnC4G8Wo4mMD3Hk0[jWfRo`c8ldP@BJ[VAX[1?0[=
GIMCWUN`FeG20U<?n=h[CEW;eGVWoFo4gMD3Hk0k0YehlTVoL4d@]lb3a[n9aH9g
Bj8C1UN`FeGZ_goS17Yl<jGDDCL9nWo4mMD3HkiVf\PS9TR4O=KCEdAf?fIb:QJV
Gqf3QnL549@ECc0lPJVQKC=M4jc3iTJfn^j^inD8AlbA=4cgST`;f?D>8n]mb1Ee
dZf;GA\T0FkXXi1<A_3GVTmkKC5`P0IQBEIYnET5bUZ>1]dg95`;f?T>86]mb1Ee
dZf;GA\T0Fk6VjjgBJFnMg;TIMdGPO>?3]cJXQD8AlbA=4cC5\hGJ=6RLV^H_S[b
oQCYK\TI]QA9iT0lj2D\TQMS=Rdhi0Mk;Uj^SH2a[CB`^jQ@>UhGJ=AI>kbmZb\3
S06bnhd:4d\9j6abjT:\2\GM4\K1T>K^0<_giQD8AlbA=4M@]cj_UJDS`DiNjBd@
DeA6L4>A7p5TJ2RkdlK3PUiG5=T;<hbh@LL736F@_@4159ZYVYFC=k836EQdPMK3
B]B[f2m>IFf8Mm<fekQM8Ol4;UBZmggK7J1^i7TXK1Gl8M[CPm>d[@`7l00D9d]6
U:44I\7lLjD5@iYe6O64a:D17;1cmMgK7J1^i706k3aNSX1`A3WZ_n83H=LM\[:7
NN_<9^TVJFJObGm9daK^aC8SIVZI3>mVFCgF;Pffk=@LjmZdP^52X[6hAQSEVmQ=
9>V[9ATV\^0E@7BfHmQ3PUimIcUT:WI7=jjk1gZ\U>DL^U5Vhc52S55n9\BQoPT=
F2d<9^75;kD5@iYeKKK3PUiGFoc5@R07@57Q>Y;:JOTmBo>EJdd;q1i@6XLn221@
3ldME[0Ho8IckhXfFEC4oWHaa2U_g0QdLhE^JdUmAJMQ^E[fjdo4L1IYWH0[]5id
JU=K8S0[<_]h=2IRJ[gO5dXeAieZQdGdYh<c4FL7Y>^InfPoF5MRlih>iC0^;5Td
J>YFi<8R_6`YAGVlo8C<lXXeVieZQBA9ShHjkYhJabVO`Um[_fC5iESAm1Ln^21@
3ldME[bKI0U^a<kfK`QBSEIMhd@\nRHFN7GCBYe?IeoNn6lMD\GIN4Y6J7LnF21@
3ldjE^GPj6:^ViI7BWk<1:@ZjWOKoA`][YSEU0gJWfM9JTLn:fC5iEL6JFJ2nJah
WQ2ViRU<WS43G0hXXpRPW5DG2@`2YnNggOob>ekf>58_gep\lQde8UbGPO]0\NP^
E@bBmajonPB5=J2\<CniebDc44]4`]TmG4fb^E>Iof:n88`O4@Ua^\`Z=jCICcR;
\Q[]6INkWkT5[51PKlZFebDc4on4e=LKaR`h;U@lbDig4ZTCY7@I^B\c\\SK<:c3
Ski3KI:1Il;BRdY;1<lmf6[Gj3QKi=JOMPRg;4m6:JOcR5R]CTZ^_BCGPO]0\NP^
NZaH1HS_V?f^g;oA[<<5FlJ`SoQ4IK@23iTLgP3W]MZSV\Ta495[^\4Z=jCK\NP^
d0]AYCS>Z2f\dnmA[<<jEWe38P63CaQ2f1W^^4QW]MZSVXCWLbPDkIce5[]og2qg
F?cL64[Da_gh@2?S:PXQmRCn^Mg?IOM[_]mk?67\nd@JVH4X9[l[5\3j<IUD`?o7
JE5D;;CCHXmFZ7Xi<]c2gK32;gP?In:W_J=KL`d\5^`N78;B<:dggB:9ZI[8`@@9
2>mbo>Mj6fed3RdUf7PBF[JnZJ_9IodK>INkGT7;^D`jdmb?Rb?gTiE9VU[g2=Qj
J=cCIe8Da_gh@2?0`Cb?YbCA7_CVdcUO=N;_V7=N?_NY7g[2aYRc[<PM13o9_@V3
F=]@OH@CS?]=;2g0`Cb?YbCA5P6X6?hagTFE^iF=M5HVB`J7997E>g5LEn@cOKOj
UB:YPHQIOeN@;o0KSoW?YbC@EE@2T?=3kUj<Tk6[]?3Ca[]kSScB4FmI=[WCLMpd
8[ZmV\dGjHc1L_gZA3U[L=E?dmha`BU]h`7IcA;3@A4mhGTBa3B0=BRZ[C[G1fZ`
I]bSoddMRea?16a>kTl6DYFOmfkj7A<HFUOe1:F8hhKUDHFZFT==WBRj[CbG1fZ`
;nnS<[jMfJ?`F;2>kZ]CdF=nYX2D[nh^d=:VcdGe@A^mhGTBa3B0WPRjHABVfeO3
8\>inSO3jH81LegjC0oUV?cm:IFU[W4^_LJ;^dS37Cg_kj]AfdPniYXC[][3^KUX
;DCSJ\eM2OkEJXBSh@JD3?amiK@FOOYJ2bLgKU<YjHiacWf_fiNng840c^4UAoD3
XH^PP\BGjHcF<Z5Sh@JD36lfE2_i0MAnE7N8<Wpoi2RC>V1jnflI[eCOeNj[giia
OCG63GBkoAAV:TLfh]NLH_2`c\a7;BhP2IR2A72S@T`:T_De_kjWP`AKM=DnoI=h
UM\V3B3Xo>S0fl1I5>XVIoCoW`AJZOg[g40b6oW[=TY:T_D<_c^>P2PKN=cnoI=h
UNRh<jkXo>S0fl1In>ESYRjDh`RU4=_EOaZF2mcS@T``\dE`U1_RZN>g:=KXUJcT
TA@@T`KOF6C5fV508;[KoTIoW`AJZOg[SI]ZNoNO<liH6hWjnT==Zg^MeSnhg[g1
TAd@T`KOFO`?8BoCh;N^KO=ahgIJ0gh8I1FeG0=aT91FF_b`BEY3AcUKLjLX:[O@
M0]Ro\SH?feU7F:<^oQ;_@kp3gf`0;@FnB`Y84?:D7@??m?0ZHhnBDB72CZ\V`0U
i0dT:DBiY=\WJlfMIWDCVli0iJI=cjTWVN?7]A?Yh@fZZdkEMHh_P83beCl0eG0<
gD7_R7mTdY\8JlfMIWDCVg;bY\I9<QiInB`Y8g:9<H@d?m?0ZfO>XD;<Q;n>i];;
m6\DYFg_M`XTj@6Xf=95l4ND3^dD^gbJTB`c]nfNgaS0P:Di@fZ^eC0JLcKQVF?C
A\NiR630SkD9j>HLVJ2\V482HgHJ<4@5nB`Y]nNU^H@0?m?0Z2lD393XeNJRmM0U
jeeBX84cbf_fcV@SeJ[@3M5Se<I_TR@NnBZZk:fPgaS0P;8faf3V\jfP`cKeVF?C
ANRRN;QO9kR2kl@MeVTHVg5_Y\I9<QiIhe3ndQ_7Sb25?8c2qRnZ22g;ZkGcb_T[
6NKJAi<nkI3]HBiRUTJVeGZOQOWI_`OP32oQ\o`SSBK@f@0jfH?SXGD:k7JGi_X4
6SFIb@07]J3]T9FoDI_<FKKO6MX>cYCEa2oQ\o`SSB_JlI@J;H7D<dK;_kGcb_X4
6]>eY27c1=fCSBi8nL<K7K:@ae9>gJ2S@\\KiD9[N?4NoF0lPR05=7BPLJ_c2_]2
>A>JOi<nkIoJXDl^_F:<kG2fbaWId<kCCW@SLNU@R<K2OmDWS@\l>[K;_kGcb_X4
6]>?;:Rndgim\Jb^fDGBhNKC`Wh>A@P8c;b7Hil[L?[\3<C__f7WC_?;kk^TShF5
db>A9]3J;llRa8UJ0D:<mG2fb?ieVYFoE\@RSEl[O?4NoEo_kV@WMG3R@?2nc;Xd
SPHBY2WI\qB:Y>Sg8I^A_UX4j[E8F^do3d^k0?n[76GPcCH:ACTaTnc]gYHUBD9h
HHA?MMn[9_3hg<FOA\^A_UXCZ=PabgAnPG^kj?PG[_R1HRFg@kSLbDLRg<9UBDWg
coUW>2CBZCBMhRV6UfhYjMeTZ_0Wh=?UNg388D1EG=5U<LHEDJHC`=bYY1hFn<\a
a>27mTVLYG\XIWjaT]52_@XCZ=MabgAnPG^kj?PGbNR1HR<K@kSLbDLRg<b6Bo9g
cUUW>2CBZCBMYKi?j9A6jDfgghYah`?UNg388D1BVOR1HR<W8;4Q]6E7[8lGKh__
ekAbgH8g4b@e3OTN8Y^A?0eNQZ:9F2Q;S3SALjh\@Dj9VR8O1p;co9\o]PfT6bnc
Znd?dUj;VI^3M^KACpFoVF?N3_KVYORAocB]41P0?X_C@AS>cbkR[:iXG:0\Lj7k
KTaZJ;CTg>9hX9X^6RMS>hVg3miChRL^R6NH\ZQ@i?_CS3M8HnhicQ5XYOeFFTXP
6k6IJ;l>Fhh6F\LJKW9cDhhOEDi`<TR^RP1W]^DL0I5hNeMYThhdi;<A9IB8e^JP
hg=K1X56^bIlC9AHX?eVJbO=mOKChRL^R6NH\ZGLB4;ULo1M[:H4;WhW:cn\L27S
\Z\IJK5XgXg=0>X6aJlS>2V03PKVYOE:S2`]59Q@mW;ULoSdj1hdi;<A9Ik7P_ZO
8GdYFGCXFoIhC9AHX?eVLc7Y@J01\LjWb8@;3qN3SZEI1@UfL<ARIg@;NXHbZZG>
8kYDQ5VFHd?FZN?P0U:D^>ofe`And_K5o0S=m9N8N<ET2bDid2lNi9j[fLH<0QH<
M8fYQB0FHFHD970W6]@nX_j:SM8CK_a3A<2h:5i@[4E4NdZEo770Oi:V24HT[PO`
CdGnOdI;XbDkmPe<Qd^[9IjgXMA>d1K5o0S=29i7:5L4c_E2RL05O2X>BP>GU?G>
8kYn1OA<SD;P\<oF?oP9;]ofe`8:WD2YX54_?Q1O\a]\2LDid2mn7JkY^1HT[PO`
CdG^Y6E5MYQ>aRN_QC^[9Ijg8KU@\TCh1h2h:5i@14]ET2G^oJJ_a`UDMR]WCiVX
I^gapIMLhD^WY70F:e_TAL<NghDgCcd>DLhOo4`JWBSoB<9622T;;63db\gR5>@n
7nSYS0GX8]@\VU]4SecTIL<NghD1C[LiWMDj<bl[bIo<gMb7_2kfBa0l<Mh?U:SB
>9Sg1IF=@OJCiId@W;caNoIX\KV1VQfHF=4RX_C1CTBSiMb7_2Am7YMe96cZ?>j?
`N7ImhGX3]@CVU]?77RZZL75;cV1V@fHS?4Rd_C1CTBj]LU7_2kCBI=ZEE<Y3ED1
19ALE[>hQ<BXRD<f6@Y5E1BFF9:<UV790R:PhAi[QnbdA<b7^2kCBI=ZEE<Y3aP=
J:ebBO74\DOLJo2Pk6IFD^5DqSckQ?__P?W2Ue9icl7XRI2V79?=6DMhRJ<lG8D:
>M`gfeRo>Oo7IC>KGKN[?;A<I^E:T[`?1`94<9_R2UfNNcVW4k;`9Ro4M7`:J?4E
I>LjVG7n4GDlECn1]Fc:lh8[9=ln`Wi_O?nHV\8RQMVjNa=iAAIo_DMhRJ<lG8D:
>M`gfeRo>Oo7IP@eCmC_8;4[ESZn`Wi_O?WiiZEXo6KNocVW4k[iQSk]R3S1b]EE
AEDc72\<nQ>JQmn1\FicJAe`cU:2CeAQ?i21@ZEXo@kX`HM7MAG`HRoLMRcV853K
jXZ]N7\>NILT_?f=Za;F2bXB:;UKq^Kb;6]bhdB^WL37bN=4SEUE5]D4cB?;`@^U
Ido<GW[SQ5C5QIDG=X[3oFZDX5[I_DX51^I@8IlfhL8B]4_hJZ8[5\]?;HLX6\57
Ae_i10TLK]<7X?KDMM6S3kgK374fNY4XAhhbjdBMWSCDJVLAO2nM0?L4QB?;`@^U
Ido<GW[SQ5C5QIDL=XILYS]ZFnFVm^4oBhhbjdBMWS4FHPPRO1nH<5?K`P6XR\57
Ae_i1a`7MkOW\ckV>k6S3kgK374fN`YX_J>UAjlDjl4BQ4YFS2`:e5ij1A6XV\57
Ae_i1jU^k=OaTnWIGPeK;[^\mal\:2LJq=<1lL>FjOO>63Q9^b?;\;ke>GMQ]@96
EMFYZJo5VaDm8DLfbW3:oFSldbFLJ@h;]UK`HjjIjXT9ZL>fM1W?I_52CIJ9^347
97219J@8hE>UnmI71EBE2V3=okFEnWcQlS1CYRiFGaT9VL>fM1W@I5FDm;3^O796
EMFYZJo5VaDm8DLfbW3:oFSDTR4kQc_YibRZeViF_aT9VL>S_\NHOkN9N;nHA347
9[QjL\77;e<UTmI71777?_8U8m[iccDiMS1O7mj7BlH>lX>fM1WIKK52nI`W:RnR
1O5jL@Yf4E>2X;\jYP]SMaM=akFEnWcQlK866^j]o1SF9>faUZ4g2oLUhi>Ypmm9
SJ\[`1K4K:UhGjP`6hcc_L9CEf851cnH`=P5KUidSI3F5W0LWSa=mPFm:6hRW_[0
Xl<[g^j_PMQDUT2FJM@DI:L;Hbfl828b2M6c^MSEk6cK0oWkZ\7`OZP;9Wc86149
8>N[U^j_PMQDU0@FSMlBKI>iC9GoEcnH`=P5KUidSI3F5W0LWSOOao=l>4h5MH6=
S>N[U^j_PMQ7H@i<9nIP0BDh?bfO8]WkKD:496SEZ6cK0o0cL@3;]iPZ029Yc14l
oV2n[[L4NYID:0P_@n6e0I>iC9GoE28b2M6c^MSEk_i5Hb_2a@H4;ZP;9Wc86C^>
GK2OL4le@O1SP[?=M3BDaha<pV109`[g^8k?:P38;kin=G>R1ihWDa]CfI6H\mnY
K4D[2j^d^0B3Ak8hdkUDKZZFCd=WO8AkSb3fMfdh3;NPj:GjAi`LEijClVUH[cm:
UeU?`gaGVdgKW^YAFD_kMbeRQ4lI_I0g[U3e8S`4A;NPj:GjAA1LeijClVU;2Dem
YIEoSj^d^0B3Ak8hdkUDKZ>f`F=ioTRS<FL7Y>EPdEKXDOTm4O`jHijClVUV2O?S
IhEO05J2Q]gK0W<^]lm^[8l464lI_IZgC8k?:LdU0E5o3UGjH7\B:D]hBaV_k=mY
@?EO:S^C572:`cYAk9W^geffBlSIUI0g[8k?:LdU0E5o3UGjH7\B:D]hBaV_k=m:
@eU?`g>2d<6YQd:aBeoNg?4A:34Zij1Wepb^47>cOCJQRVoKHmHZL4CPY=1<[HKD
cU7Tn\k=2RA909<a??V[^SbG4;fFbjN8>mNZ^7>gEaL_VeN3m;Bg^GQ1nQ1;`XZT
49JB4bhb1NCkQV2am[HSjcPJ[bHiZ4V6^CUB6a2amNjbhODd_7Bg^GQ1HEA;`DZT
49JBEbHTl]IG@ZQa??V[^SbG4;dH672A4O0;4\?MoFGa:TEgi5eWIkJRLU?AD4ZT
49JB8bHT8bAjM=5OSDQSjcAiiI4Hc0HJdIUBdae^c9OQ>GNK9d>g^F?6QA4fj=G0
S2JBEbfb1Fdj7]6ngE0aLIEJ[6Hi3kQAY7g?=7^eOUJQRV[LOMnW?k\1HeV[jNn^
BgZDkVfb1FCkQV2MSGc2W4Bfi0?@?554QjJ_BWBl2;qT6Xj6Y82@@Q?CVf??<n?n
P[[ZifI@eJHBR[Ppcb5GOFR2:hBo2?U@bXoMTTfN6:ABTTMhWR\W0ORVVKfKHUB:
Qf?]2Qfi;_j=k9:0_Q[0[9\HgeL[@\ojh1IXh:Tk75YRB1APf>\On7I6Y^[6T[B>
>c]=^YG`5MNe>:c?<PfS[9\Hg8K3@\ojh1IXh:Tk@[IggTZD^o=ji;gkIK>?GK24
>iik4<ROS:FJg=ek<ofkBBZJ6c@ij5_MAOIUh:Tk61a\E88^VRUdR6IIYfo3Gee9
>GIj_YGRnk7a[mI<F6a1M9\gG[@GCK<53AIOh:Tk@[@CBG8:Scoh5OY4>B[UTdM7
>@RV0Q9OST2m4c:nCGao3VZlIBK<@Rni54N9_:4`Z[@1B1APf>l<RITD;N[HbXN?
4ViJ7]n>n;^@LCq@f2S7mA^Mh=Tf=go_aKCjg`6=jRTb3gjDoITm]eIZd1o[cmJ3
Rj^<_Id81H:\akd6^Q?aL2YJaN0>b=@FiZ`DB=II\oQEDnf3;A1NBCbJ2]kIB[Om
KEkjTBQTO9SBj\HhMXXHDWoZ`NA>3gQLWgM@B=@I\mQQ=nj9YfUE=ZMN7]k5an31
=9@h7RNhV3J2b4BhjG=bn<;Sg=Hf=go_aKCjg0FoD5G1@chZL;4ROZ6N7]kIB[O>
KiKP7MI<CU?Y`iah2PbbZ8<J`Nd>b=@FiZ`DB=II>Fo8BWAd`Cg6]Z<N@jS1PUKU
=X9CF\N=YAkH1kWYMPXR;2hjkCH:\=a?IU9:B=@I\mQQ=djZ`Y<E]<k:WgjE\OJV
oTN@^^ZFVqlXO64Zf[:eE7Wo9FKk3F:MS^A>58ZMF2WL]l1nLC^MdH5;i2\8_bAe
8<OeXaJ@O7i3oYC3]K:PgWU6WnI62?AV^a@Vf9o3j;C88G?jnNUN8oT5dUB_YCPP
h?2P;[@SHN;`e1LgZPTeTL:C]DI62?AV^a@Vf9o2jFFD\6Y7QR>MJg[DjK6UCAgZ
8Jd>=dZBUR;NeKLgZPTeELWo9FKk3F:OSgII7JW5Ui_X8Z>lQR>MJgc^f6B\CGgZ
8Jd>BKiK<Mi3HQRg`UP4ImgjWWI62?AV^aI6k@CBBADHLU@7QC>MJg[DjKIUf6@Y
87n9_CbK<Mi3oYC3APTja5X6287G@hDZA1MkojcDYak0p3Blk`YcmLijH2KhM1cU
Ii?Yl0N?bee_]<=BkFI\mW3`jXNO<Fbo^X;Z642Y7Hb]3f5<G`>cH4[m=a9KYLSP
Z5fgnJKBnAE@i[Y1?nILM5Y4G:0b4\oNLNghHG8^5G>SB<8H0UEPK7`m;a9KYLSP
Z5fgnJKBnAE@i[Y1?nILM=@iSTIcVXDXK4SZ\imSKG]G^<;YQUb\BAWAQ?Khn1cU
Ii?[G?XO1d\CRiCM<LJL2=@iSTIcV_mMUQ6[TL>1<07DCf5<G`fQ@4[m=a9KYLSP
Z5fTO[aG0i\`nZCnnWfZ6T]mm;LONnCqFP:^d_<0i`Am^:e_E]0SW;9Q:@9Heod[
o`HgI:5KbF3f:I=DiogDK?W@LLA^K_O]c?;YROPYP\6[WZ8BZ?@GK6<KchQd>=h4
=2;FYIh;_UgiMl`ijDIO^Y<SZZhiNUZbTdEm[kPJP\6[WZ8BZ?@GK6<KchQd>=h4
=2;FYIh;_U[F@X6F14IUAOWFGd\W]ZDV:kNIOiPfiWVX8^nY_0c\W;9Q=2]5?dLO
=UJ05Ohl_U[F@X6FUg02W1T2ijOPkC[;c?;YRDOHP\6[WZ8BZ?@GK6P9g[6Y6d]G
]NMAdHb_>^E968efmOplj@NMgVki4J_Zbmc:@=b2]NLH44ni_>3oI@ihBZdi]iPG
[=\6HSPbiQ8=LAW@Vd@80S[^9:kLJRC[c3BV0K=YZPG?aW07C]89D9T:8MKb\cTg
ReTiJO8GjFE?d_JebY380S[J0:YLJRC[c3BV0K=YZPG?aW0?R7J`5@C;:Km2;i8G
[=\6HSPniQf=LAW@Vd@?5HIh@MX9CFo2=nJm8K3YZPG?aW07C]89D9T:8MKb\cTg
ReTiJO8GjFE?d_JebY380WB?2VRjCZS\ajY_6h\^lZ<i;F_\mqL?G@G>8GHFQ6J]
KDPg\@6OJOCjXl\7]BOo]Bi3@Uljoo:6><ZE3YoU4`HR=mh]HD38HKOXo=1`IlJB
2e]h@76L=FOme4F2OAJoK32Yde3^A1m^S9ffiani3L^kK7UfoD38HK5Xo=1`IlJB
2e]h@76L=FOme45JT_Fca6OT@Tljoo:6><ZE3YIHc8;f=okOi3g_1T@^lN\I`o7_
OOjh@76L=FOme4F2<IZglC``N0ZjoUm^^9M_c^KHJ]9kK7UfoD38HK5Xo=1`IlJB
2e]h@76L=FS]BXEPRLZP:_DR]Re5emTNS61i]qN3=JNK0hMc\<QZlUl9:3ggF[R2
lnAS7<;O8^aQdUR6G:I5LnQB\]>YJ3iQ>jd2m8:H]NSbo[Mci:O>dOc]CTaRhA18
AThKM91=VcRAK8W?NTkd`9>3Q0:n;LhfSnBLh0?9<iMcC<1QZPO>dOc]CTaRhA18
AThKM91=VcRABoR=D[d1:8QB\]>02]]HACX2?X:OM0AMJFhaQ<^NKGlNZ@lS_kih
66hKM91=VcR8BkR;@^djL^OC1Ma?XF1B>:?2MRXK]N5GkWA`f66QLklgiB2RfidI
ACDm=O]OmjhVK8WXEgkd`9>3Q0:n;LjkBOAOLBh4hbI_ihoPQ_>L`6N0Ep3^R>Xm
18<DTYdcT<hIBoO@AQ]ZU5jSTAP_BYnj7Och?D;gZBeDfMZ_iYK?>BklnZAKW90b
lJjDo;hF6m4O5\>d>fb6o`G=DOA3N>TD2\gg1A;X88O?f_>OkW5nhjI829SEPoHh
1C4odRhF6m4O5\>d>fb6o`]dZYTml7^h^Ym5c_6J<RS3FEoITTJ0c8b1nP;4Z2bf
iZ=:I]ZWZ`f9mR`b0eXlo4G=DOA3N>l:T3F5c<6J<Ra?DIZ_\3TSD0hl<ioRa`7h
6h=[_?A_T<fK=K>d>fb6o`G=DOA3Vnn\_@Uocd@0ebN^[U9eAO1=IOScqJof4[6h
jA2mT6kHVj6:f7XJOEQa=_=k?3n8AJEEQ<CJCqFAQ`a?FVB_j0hT\X9MBYSVPS>2
LoLo5K7=HC>TA5iXjYHVHe2mCA7JiTCY8Af=_Z>d3X]H6IZcjK=0Q_G]HlWlO;8i
KS38IL13Y?bBe9hCU7ho:Zb:W>kIAakh4oOAiclAJ>^_FVl[gm@0Q8G@5PSVS?7L
G0\B?ALV2Y4VNnhCU7ho:Z<mV]nfiEZN4LOkgZkVW6]NkVFCf@mGI>5b^<5=G\5R
3R^03FO[YhbBe9hCU7hVZcNh9X7fTFPH2\f=hCjiOW29B7WLYJ:2@756^>ZVgd@X
3;<HIY13Y?bBe9hCU7IY\::8g`a1X]LeW[`DGO\oVJ8f0pd;UO=lS24MYjg>R;BA
UVc<eD5AZ=ban`j8GE;:OG\E3Ag5EI]SMS5KJdlGI>a=KOTG7Igj]4nEO:o2N=\B
9gI0RJ7S13<hNnh4K9LLW\?FR@RhI;g6m9kYHFR5[[lGO`FCgXGSS74>TlNC5WE>
S0f8JYQ:Ml[hNkh>nHMLWM\`BDLiHgmU?B3Ko6@fYEbBI_4D^DGSS7aMY0CTR`A[
c7W1P?UHZ2JdQFTdM;_akEX43>RhI;g6m9kY_iZ>glocIM]c^S@9Uj>APZmACJQ^
lZND0=UA:2@dQELdM;_akE?FR@RhI;g6m9kcg=BZhXcGGPD1`V4mEEEF2H]_1JpA
E:HZiW1DkkjcDPeZ6C=ZO?aH\IgfNlE4dT]J^oF59HFNiX91=bjZT78L_YCZJWS7
a1432ic;o3Y`5R17L0B?@^KNF@K^9bojXEhLCGJP]Ko^j3H3@h`_J5:n^5TS=Y>E
`6S3`WZDkcYC;c?QARh=[=?KF?5RHiQ^4]In6MKkc3gJJ1A6h8XLJ5kn^5TAXVT?
KL=12jAP_h21IWlOS<M=LhgNF@KRHiQ^4]In]aEI@VBZ?6PYhCf2]@<XPff;0OS?
c8:NAdIDkcYC2W1OL0B?H_c?ilm44]QdYAZT6^QN[cm88TAUJLfCa@>?PfaR0Oc?
c8:3`WZDkcYC2W1OLJ^Tb`R^9gMCfL5X7ff]G<=;EkfPYpC79ChiMNlj:EFK@jXH
H81P=h9M@J3>nhMHT=fUDcE6PPPA9Al\igMZ^_6l4iII=2LZ^>aoTD_R^Jb>5TIj
;mO<=DCdb12N2K\Ede`Z`dbKGWTY;iZE8WYN<2A7o^DjI8LJle_FMXljch]ScnOn
HH`084CdP1:oEhafGO:RU5Q8=CSeA:ISd=lN<gA7o^DjI8LJle_FMX_jhWKic4On
HH`0849ME31i2A\Ede`Z`dbKGWTY;iOnT5R0^jj47e?g8dC`EV<VchOBM:LFKFnV
jEZW2BINbo2N2K\Ede`Z`dbK=WYeA<ISd=lKQA0R9g[ofmgD=TLhqOPYX9;<h9\7
^[fLYc?X0VXDD\b_lYbU^9=RM[DRAH75@OX0AYI;`S0LQ:j\ELEUlSYIXbYOPPZ5
a_HA>[@X=\3aP726g>iV@G[BHLUeb:TFb\]MJo14RjZ2^M<fLfUkJe@JaMB<k9\f
^AfLh[@X=\3Qa726gWP=^kJ1VBUm::7:RSG]b2?]mjZ2^M<fLfUkJe@JaMB<k9oG
DLHfM0n>BjmTlA`f:F9n4LOBI=k?M5d4SRn7bfK7BVZ2CM<fLfUkJe@JaMBGe0[5
;hHLjG?2RjJJb01:Smb>N9AFS9F7hlJed\]MJo14RjZ2^M<fLfU337:8O=kF_M\U
oRGWR8V:TEWL\?dqWg?[D5@oNSS9L;4ViC]Ko_3:6H?8FFCL2;mNX8h?mgk>ob_U
mLAeDhk?Xc1_Q=Vn74^\m?F\Enj6:CX0H`G4N<BR5lh2=B_h98G73FN7aR@5_U_]
`:ZD<l9^l56ZL=:8nacI>6@kNSS9L;AGl`GTJJJa`=eD\;MF]gLi?BTJJ_a__Qa`
m:We?XkeXc1_Q=Vn74^\?aBT2734]oAMl`GT:HlDJIJVRM=be=50;191ATHOdb\[
ALHM8@4Mm56ZWm?bmCc;jN<_`GX[:;AGl`GTN<9?RgST0RKb][]mIF=\^W@HI8VO
QAQQ_bh[bg]]XL:HnacI>6@kNSS9L;AGl`GT:H[jRIh41f]a5LZmUF>T=f8T=0ep
d`=jIoP60XTDm7>`YKH9EfhfdE;o:9>:^AqYYbkd>A8\6Q\Z8f;bXPN8EMWCZ>Yg
;QI`4ADODZXCmIW<GJOG\301NBM3\nPZD\FkN0kiPeePINUmLjfnU;YBPMO[6P\d
]`i6JABIh3KU[eEX6idgYGm1W0J<AE^n8U^Y;<NDOAD\6Q\Z8f;?@RKHjj4iZaid
LBAU;0JIh3KULEE31JNFf>S;oBQ3\nPZD\FkN0kiP>1W89I^ndE0cRJ6<KMhQ<L6
UBo4TVF7Tn11RDfdSJJGh3^OaA@Zh\iC[HN?;<fDOAD\6Q\64_6RdQ;NUKMh88i0
loJ>IHiIh3KU[eEX6idg0JA1T9SjO\\C[HN@jh^FC:;EdS]2diBPe5G\8;MO8fpm
LZ9P[<Km;:fiI\o]:mad[B?52gR96To6<3WjX;XN90Z3W6=\kfN[YT[1mQYEiLXl
Q?UVECDjGcRlP2LLCIg2O?^W22UMFTK_8cIJ]S4N?[[F83oQ3\o\KVLR30TEJ?oG
i2_O5@<^nePVP\]]:c<\HQ_PTML2jT46<\nIBbci]Ya01<JM^\`NONQCmIiLiLZl
Q?UVECDjGcRlP2L`X8:dGB052gR96T\_8cIJ]N45][XF83oQMUC\ZNeRKm;?8CLd
>n>4M<Rm;:fiI\o]:c<\HQ_PTML2jT4_8cIJ]UQ>V=7U1<ZM^\`e6_7LZme>BEV3
NO4f97:X7`\X^h1pAA6P>k<]l9B3[cTR?J^X:3@V^hno\bRW<`OmnnBjn@Tl6<fD
NCD0G3^[2J^oJ@ePb=TiZVfQ:MUcbM1HJ<_lK=aYTUcEV\dQ3IMAE2PenUOWo9Gk
1_W9FFG]Im@[VKe:WN0TJAccWPFHQXTR?J^X:3LdCUeRajdV``O7[WP>nUOWo1]7
1`VNFa892J^oJ@ePb=TiZVfQ:MUcbMkV\jacY_fHTSBJfjdW3IiGB^J\3kWDI\KX
Qdjh_FT>7IS2oCmV7cmYA0;=l9B3[cTR?J^X:3LdCUeRajdV3IiGfoGeQi\<Q@]N
1`VNFa89Y`^Ho5>6^BjVo5Fo3@gPXFa:qb4g?9]Rj[i^[^RccH:m6[mZ?bSES1a<
?49QB>9nDVDlmLX[K4c;aTMXc5<R>f681BbX=@ULK[Ph`Gb09lVG4a5g695^k<F>
^kfLKCaf83mZd2c[ZlC]7TCg`GMQ35l7bQQ5LHaoQk_R[XL0bH:m6[mZ?b2Z1]F>
Ok]2Kg0[J5WbHPa[GlC][SCYV]YCNf^1H7QT>@ULK[Ph`GbH_L17HjPgC9;G<]F>
OkY?[N0[G5WbHPa7R@PZ@TiVLWO^L@^]Q0ghRE<jf[i^Y^RccH:m6[mZ?b2Z1]F>
OkY?[V;V;m6f>`cdYlC][SRjV4VSPfMPN<MknUKKl^1F7Va;mpD6nD<EFXh6F\A^
6RMS>hV03PKn_;nfmiEZJBkX6WPBmhB7@TLm:PPDa9l[5;db;nG^2ko0fdcjAI6Y
G59c@jm_VP[GW[DQ[:E_eV2Xm2;UX0E2S=L0b0@g1Vk7SSZ580YB2UCOfbF6]RfY
Zk=c@Nm_VPRBY:E:S2`]59Q@mW;HY]4R5=]JlWnfRAoYaJZ580dYFGCXFoh6F\A^
6RMS>hV0[fKPW61fmFEZJBkXL?3HY4><k:mjlj]dI7oF]3iDR=dYFGCXFoh6F\A^
6RMS>hV03PKVYOE:S2`]59Q@mW;ULoViYNl00lnDj3NURZQS9]Mdob[Dnq[Ed\hX
a@06dMDB=;X<iZ@jn^K^N?ZMZZCY^\mlY?A]kSR?_PBLeooYEZRH@U\FDE[XbcnA
]GkEEYSWPZcM]7_n32Kj>CJW7P4bMM]iF0^YY4U5CX:ig7gYafGDFC47]Ujjhk7L
K3e3S[P6nYX<iZ@jC93\CkJf=JEY^T3S5@l>o_Rn[b[;^iAoEJGAFhDEXCTfc\TL
=nP8]=LZiPl^OakIOCho4_o8oC=HWD30bS_hG`WBgh7dF[T1alGDFCDEXCTfc\TL
an06dMDB=;X<iZ@jC93\CkJW7P;SQ;R8FE__gAMmLY2R0456TKf05Eq^1;b<4To8
`4ML`TKX;KmalcWYNKi]nEQbN]f]_FlAAj>>?7acUTQd1_74h:L;8?_k[80DG;UE
D0;6:nC^J>_KKRMdb4hQS@nTRleWPio5MUjY^KLO11B\4^lKKNXGek1<[VGWhij5
\>S6VSBlZgR27EEU[KnLMJXgW>>EVX@\;=[fI`YnhT@km0=jW;U[9X@eGQ\@b\?W
\1[mGCecF6>lBg<0YXn7_jHc@=5]kFT?MG;S<8:O>TGjAm5aKN`9VMeNlg1M5T`8
`4ML`TKX;Km=NoC?8^0HJMU@W>1EVX@\;eGP`l4ODM9;Ke529J;[RYCLfEB[2qJQ
c@D23L[YY6\L_LREI`IOCHTGZPXU=f?CW7XRecK@@nMC5SGRAD^`D>EKE:[O1g<6
FA^n?>NEn5W2aORR=9U6NUlkgf0h;W9lGJ[68_9I`UbGIOC:b\FR_Y_7Z0SibUJP
fmN_U_3:LA_0MG[Nm@R@DEJ6SIN1glF9CR<I8F9DDmMc:l4J3ZTUTOFG8E[LSka1
meN_U_3:Z[R2H>4cF^KkMilH04R_=[\T_bX65ODf[R1P<afNZCJ>F^WRHgb[L[3a
58VE3D[YY6\L_LREI`5Z_AD6S9N1glF9CRb9OG<9[mcjeQ>Q>`1Zj563>V8TWqOD
j`;S=oH_?^Bh9ZUK7bD6S5YAL65=OZfNdTE@C15Vo2<@Q=8o89SY6LqEAUTOO:U9
1bkQ?RgM8^@3jFfbMRTmkk6Vc`oSQI^:o7:foQF5=3?P4gDV@dPi=Gg>j<<`KijS
22?5^==GRQb5Khb]eMZMkk;V>L5mT>WeOheKl`\Y7JlP\Ml:ULdi09_Y6EPO<0]i
A4Q?7P>JE>jRVd:`O<:D@NcoT=GV29;PIR5\bD0F_3`64R1md=M7>bFH3no0<lXL
M=CdBC`DM7cg:i2YiielKkAI28QS5>fnn2QhC15MlACXD^Ok_J:D\@\6NaWVh:L9
1bkQ?RgMcJ`3CUR`O<:D@Ncokhla8\:6N2Oekg^>S?[TDZ5k6_[j`Eq=O=]K2?5d
44Ra867XU5]ABZB<HYg>8@W36d2n0fAaCS=Umc\FPG][HQ78>Gh6o4NFEYnhHG9T
Eb[j2@0_U^;[7HQ=h`[jN73F?eKGglLZ;6BEO39>jlhWWZQj>eHfe^^^nae^\FhW
M58N9][o]PC>kH@fg_YjUY[3g\\Kaf0F=P5ELPIFjeHLHQTQ4QSE<]OF>G9J2?aK
44`aU64CFPj8XMi<hSOVPH68g;Dndf\I?a\[330GG6YC6B<EfL2`h\j@iKkA[PbC
E`<eIm0_FA980QQgh_MR;@d;e0<`=NkH7@dcd2]\d>HbN3lj@:G`45clcJjYN?Xd
44Ra867XkfiXDMP<hSOVFQU=KD>6`YL1>OBhQq7U:1mYF6DHi]XN@d5=UL^=?`UD
bL4fNRDOIYK@nPTNfRG4AK3WiTS>jHkLBR8]Q>;SRU\Sc<0hh2[jk9gWNnh[d_oo
R82^W3J7;\29Z3f@RXV09A5mR??d0\kLBR8eXB=5QPKdgj02a@_N?DeimT8n7doF
W_BAWj5DIVa6PHag5SaKI=hBleUH0GO>chnQQjdT[_h]FGDhY;_[P\21m_`_EaP3
5idNm\\KIPaaIE^NO;@`9Ka;4VZaEU1^[JaHfiDbA5XX92V70N@TbQZ1^_oa?`A6
G:QXLj9g;?fT6M_CVX^C<o?lfJeZ]mo0cP_6jeUWjjBeFGDHi]XN?aeB]=8a\[J<
d5caE?S4SJP=N5XRqR6J_YGW>>oE1YR2mQ;U\2Sl^o:UW4oeGiPW`BeVk@nHVZW\
[1_27m5hXA`j1H62VA4c?=9a?Y;WQW4L7?=@k]RRo>D^b:E;_^iCj8ZRl=h4`>O1
<NUE7W>8h49UU21_B_K7751Y0M[=Lb6EdG47OWMng83J7_>]GVIoOOCQnWhdkkcm
cDA8>V;CLV[FId1AgR5^<EG1LiP5[KQ2CPK1KiZB`<MUD4o<_34<P;DZe_I0XBOC
HC5fQkEhSAoekLPfC0U[LFTmhELWRK`Om<EPH0]bW^FVT^>][VIoOOmkO2\5XYKR
\`Q6Fog7j9M]7Z]:]aYKRAaWV>oE1YRTV_PQFdOQkmFJf^>][VIoOod3md5mTS5X
>jBR5q>\3Nb133?DmRec^UnkhocXZQYE\U4NQdWTO^FA>PII@fQZ=ZXkTgf9lKA^
9^>F=gi0^NSAA6AhO0nZZNn1J\\a7fE9;\h_aSkT\eFom0F_@FmbBC\3^kbDTbLk
IcC5Qa>5Hbe\P0Cj:]RV6JUK@QkGb\K9h?4na<;jRLLk>aJD>:gc=8?XodMEF:G^
9^R>oM2@k0DOh`=7b=\:B<>XIO\a7fCoR>[H]`Ef@8>J:TYV719FB>hXW1=`coCk
INC5Qa>UU_6]3Z?DmRec=U9]FZa;c^1m][n`iQi;IX=\J>\:MS`H05Fm8MR`TFCk
INC5Qa4:jmff^V[[mcOaB;pXolgk<>AHV:an2jEEbgORQVI`dfkYJe:Pjko]_8To
92<2Ho;[5j8Y[^0G>M5V4LYlDcPRDdmdE35G:WO0e?8J4Q9V4lYo_j^PjkoVPYA9
<iIbm1kD5jMY[^0G>ShXS1XUSdBgcCW`TiD@YWfEXgLRQVI`dfkd_]QX^?:4H8Ia
cC?MgUQ:50WiFio=T81XSL1nkAnX\FV[b@4fgT8THOJc?]P:df5P<BULd1m\:CPa
9C?Bnh@\Kib73F5]3cgOZ>MXFMog0>OHV:an2Yf_AF6L@T]D8SW>8KW8V0QZ_\O4
[c7eh5gPQZ1\32h]3cgOZ>MDEg9CLMb3:bn46^=q;Tj`F06Q[mUOcTnPI9`T[]CS
cZlo<62qC\<UgnpZ[C9^@XGWGl7NHnpCa`lV[pE4@MG4O2p:_0O]O^$
`endprotected
endmodule
