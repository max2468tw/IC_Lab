//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2017 ICLAB Spring Course
//   Lab09      : Coffee Maker
//   Author     : 
//                
//
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.sv
//   Module Name : PATTERN
//   Release version : v1.0 (Release Date: May-2017)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`include "Usertype_PKG.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

`protected
cW5[QSQd5DT^<L[DF>3[glT:P9aqEGAIY<l6V=WK1WOB>iFlO0^CA5_bpcB4FccA
[\Nd\A5mDf57m>jUVS@^MBfJ:ZNnQfb`0>RISO3?]`kPWBKOG8N0aY0n=p851^n4
q5O4oAfH;HK[SZ\b26LYYGg3FCU0WId1QpU06d1]Z>cEHldl;5ZnMV_?E7YS?WOO
8AZVOLqC]hQD=JL;Wf>_Smk;dl72\5f=2M[d3Aq8bMHR_bbejiDnn4nF@\hU0GoF
XB2K3k@?U15@mq0XnoVe]N9O0o>ChGR01BbaRkq:emT[@k^kLV9c4L@MZ`T6`Al7
EO0Ho<Rp=c`^A]7C74dQAOXY8jgn8`ciV66A[cA[]WY<3F;IL_6Q3j[J;NHR?]5]
C8pdFYZRiCXa_GE;T=7m^;j8@j7nMPK]O9Koa4]?1LjSmVb7PEULe7;E\]F>Jq6F
LZMVlQTQoMlg94\TS[NNH[_c1n<HeVR8lFAZhfeaEj:gNT1?`48UA=XaqVhAfUEH
OjiDcV\8L5g5T23^;Vob=F_F>\f[HfJjWFYk_O=;M@gJ[AZL2F1qGCU?MhEUbU1[
KIXi1Tg2JNaHFddN0cDp`BfgPDPSeZ2]OV2>_@\X\6IP^0dW7<0k26gpE40ojg<p
Io^oK2_2SQkQWh11oh:ZA1@B?EpFbcULXW^ILMKFgjTbW_aoCL@MJk[@<phb=66P
nq\=P8]_mB2H^Od:Zobm0f`Edhil8WVSjf3WC09J@nJ5=q6\T`;DVH_a@Q`cW^HZ
GYCV=M@XefTJ]^nXXij6Mm2IQq5Sc4^eVoo2il1<Z8<aFYmU7Om:e]Hic<>ER2o@
X[VC2q5h1nWo]B4WnaVTBN?c8Q^77jdaI_oYE9]Lgh]aH`[f4q4c\BD6XpeU\m=n
E@odl5g^74pUnoVBb]4>@>7Pb[A^G6;N?lG4^g`>eDPee^g0Z]@@Bq0U7AXKhU=A
^53KLN@G3<Vjc?;BoUQFK^`0pOa\_2f@>m2I;;2_3fE_mFGU_VhQYQ\m9J\3WdjJ
Cq`3eBYK0jSLnVY?[VN\g36P<ccY4VjaEq3e7][BLlL`Ti2Objo0bAWC78988hE`
R8lI2q^kPTUSIqT2KGGFc\dKI1<0R5gc;PT@dn;^Lm09qIbnWS@2q]c1?<KA@;m2
U<2><]7==35j]HXSPlmgS7ELYa[MD:iiI`=gj0_e686ld`Uc2LD0pAnL3<GdLZV?
`R[aFcSVM5bVD6kA>e]PEiRfE\A4>16YC<9_djSMp@CGgQ6Lq\YPk=PM:_7;Po`_
0qYO>>08c9Z0Z\1YV5UK<S0dQCHj<;ZPmpiU^VJFU_i`==^B_YR0Ijfm5qlQRf9<
kL\DE]R8CMm7KO29ib6H>g@[h8imDqgiX\O6_3nX4WHSEVg7XY1PUUbMjS=Ddqi0
Rn8\8S<K\i0[N;;NLCOn^GaXk0=Kl:_[2q=3hK^^mqcm]K2c@H[T;B_Q5_@B@A_e
P>Fc0l7lqNTbF9JRqb68`g1Fk[K10PHLLI<nfSMibWA0G7LJJ=^R[IiU_[S^h<Nc
QAM3q6M]UffNMIUGVFSRcCApG`UNQ^LqDh[Ofog02hD8a3HYpXl5[MnU>F:lHJd3
>e>`9B7WgVHPL293hp\fEcZLTQ4]l^hnOfhcm0Gc4jn_BRjGk7Ec2mh980T8L^AD
g[qVK\ZZDg34_<O8NA1aaXclSSb<`AEbWB[_??TFU<QcZlpEAmY61lmaD31KEf;@
GmY;8g4]BVDGnb0DamE=[@oYGg2YOMao3qT\aAnYIRCGg@2eY_ZXM?Wm44<5R[1S
g0bdeC>[0JJ`4;qFMO`T<gd3\;SKRjLl`J=4F89a2AUVIgqBW:Xk;onoei3V1n1`
PcfpJ:8E`h<K=CNe7MgXiQm4AF`[Mb>d8H[4LQ;qHS7fdU]qo=RbnFV<?kdJ7DPN
[g<IMEb_C`NlH=q03`N@:TqNUFIBBXijh3X]mNmcn[8\=KkPFH5[VO_dX_H7WjHW
QkKfO3lP`Za7JIF=nHjU@AECATqCI?QXVGp1b8Jcj68Bm<9HRS@q4IlSG9]9H8gA
fS1cca8gqP^FWGXI^?FQ`Ofn=22=<]9H5V_E08C[P8>3;qM0=NReo;^8GE@Lk4kL
GGNJHbKY;0kikVF>p=Pdo9Bc1fD6cg4iLSST3idiC0\D7S9nqcUMS@PhgDhE;LGD
:mJoIdIb]VOLQ8N`<RZdT@LdW:3?Td4=FX1S5P2^oF4XARMYI\3fT<BpGjN\h737
nIg:AL5MAM=02>fb;k<M2W4MBJcqJVod3XDqF@1dWn1Jc8?;MaJRkS:^ON_<7L3P
h2plAnbF7>_H7_552WJMA<KWQPH3:8JCXhlg[0iaBf_5e?P]S8^q1YT5X=8qMY:2
HbN6?nPVAIGL;i?XVIhKTKZ<AOA=kWAfqnO4U8jHp>X@QG0PbOh?7i<F>QQ2ihAB
p:625RVC9bT[nJ1=gpXZ:m4]NA0=8>@>e][BHlQON]fBQlA\>4iAVbAG0aKE4ggN
YTb8cK106@\24oDMf;F3q6ShGW>L=Bm[[BU0Cjdnl9THI:Q1dW[fbIX5;Pi^?cPW
dYg;;1keEVGedciJh`?5b@@7DqSOFWofg]Nn_MI]lM=E2H^o64M9?Bc859U1lSCV
OmJSA@9S_;BLT]KB=OPUkOLlGpj0P1M1Z3gB=U[_8dHC>f_?5iS6M:6h>>GjmfNb
\XJPTB;iRLLPgFcn;XZR;B=D`g]VpS=Cn3FYhHoQ_6`J:kEeAB73jRHB2:d_[Ng9
^:09U`iEY;97Q?2R\80b5E<dnUoNK$
`endprotected

//---------Recorded data of CM----------------------
ingredient_window machine_info_inside;
flavor machine_flavor_out;

int supply_limit;

int i; // random initialization is successful or not
int iter_i;
int iter_j;
int iter_k;
int iter_total;

int gcd;
logic [9:0] capacity;

int check_output_times;

logic [9:0] required_espresso;
logic [9:0] required_milk;
logic [9:0] required_chocolate;
logic [9:0] required_froth;

int total_ratio;

//---------Main----------------------
initial begin
    reset();
    for (iter_total = 0; iter_total < 5; iter_total++) begin
        for (iter_i = 0; iter_i < 4; iter_i++) begin
            void'(select_flavor_rand.randomize());
            if (select_flavor_rand.flavor_in == user_define) begin
                for (iter_j = 0; iter_j < 4; iter_j++) begin
                    void'(select_size_rand.randomize());
                    for (iter_k = 0; iter_k < 200; iter_k++) begin
                        void'(select_ratio_rand.randomize());

                        input_supply(1);
                        void'(interval_rand.randomize());
                        repeat(interval_rand.interval)@(negedge clk);

                        press_buttom(select_flavor_rand,
                                     select_size_rand,
                                     select_ratio_rand);
                        void'(interval_rand.randomize());
                        repeat(interval_rand.interval)@(negedge clk);
                    end
                end
            end else begin
                for (iter_j = 0; iter_j < 4; iter_j++) begin
                    void'(select_size_rand.randomize());
                    // void'(select_ratio_rand.randomize());

                    input_supply(1);
                    void'(interval_rand.randomize());
                    repeat(interval_rand.interval)@(negedge clk);

                    press_buttom(select_flavor_rand,
                                 select_size_rand,
                                 select_ratio_rand);
                    void'(interval_rand.randomize());
                    repeat(interval_rand.interval)@(negedge clk);
                end
            end
        end
    end

    iter_i = 0;
    for (iter_i = 0; iter_i < 200; iter_i++) begin
        void'(select_flavor_rand.randomize());
        void'(select_size_rand.randomize());
        void'(select_ratio_rand.randomize());

        press_buttom(select_flavor_rand,
                     select_size_rand,
                     select_ratio_rand);
        void'(interval_rand.randomize());
        if (iter_i != 199)
            repeat(interval_rand.interval)@(negedge clk);
    end
    pass();
end

//----------------RESET-------------------
task reset(); 
begin
    $display("*************************");
    $display("****      RESET      ****");
    $display("*************************");
    inf.rst_n         <= 1;
    #10;
    inf.rst_n         <= 0;
    inf.select_i  <= none;
    inf.supply <= 10'd0;
    inf.required_size <= no_size_inf;
    inf.ratio <= 3'd0;
    inf.flavor_btn <= no_coffee;
    #10;
    if((inf.out_valid !== 0)
        || (inf.flavor_out !== no_coffee)
        || (inf.window.espresso.led !== red)
        || (inf.window.espresso.monitor !== 10'd0)
        || (inf.window.milk.led !== red)
        || (inf.window.milk.monitor !== 10'd0)
        || (inf.window.chocolate.led !== red)
        || (inf.window.chocolate.monitor !== 10'd0)
        || (inf.window.froth.led !== red)
        || (inf.window.froth.monitor !== 10'd0)
    )
    begin
	    $display("*******************************************************");
	    $display("*     		    ICLAB_FAIL      		      *");
	    $display("*output signal should be 0 after initial RESET at %3t *",$time);
	    $display("*******************************************************");
            if (inf.out_valid !== 0) 
                $display("(inf.out_valid: %d, correct: 0)",
                    inf.out_valid);
            if (inf.flavor_out !== no_coffee)
                $display("(inf.flavor_out: %d, correct: no_coffee)",
                    inf.flavor_out);

            if (inf.window.espresso.led !== red)
                $display("(inf.window.espresso.led: %d, correct: red)",
                    inf.window.espresso.led);
            if (inf.window.espresso.monitor !== 10'd0)
                $display("(inf.window.espresso.monitor: %d, correct: 0)",
                    inf.window.espresso.monitor);

            if (inf.window.milk.led !== red)
                $display("(inf.window.milk.led: %d, correct: red)",
                    inf.window.milk.led);
            if (inf.window.milk.monitor !== 10'd0)
                $display("(inf.window.milk.monitor: %d, correct: 0)",
                    inf.window.milk.monitor);

            if (inf.window.chocolate.led !== red)
                $display("(inf.window.chocolate.led: %d, correct: red)",
                    inf.window.chocolate.led);
            if (inf.window.chocolate.monitor !== 10'd0)
                $display("(inf.window.chocolate.monitor: %d, correct: 0)",
                    inf.window.chocolate.monitor);

            if (inf.window.froth.led !== red)
                $display("(inf.window.froth.led: %d, correct: red)",
                    inf.window.froth.led);
            if (inf.window.froth.monitor !== 10'd0)
                $display("(inf.window.froth.monitor: %d, correct: 0)",
                    inf.window.froth.monitor);
            fail;
    end	

    machine_info_inside.espresso.led <= red;
    machine_info_inside.espresso.monitor <= 10'd0;
    machine_info_inside.milk.led <= red;
    machine_info_inside.milk.monitor <= 10'd0;
    machine_info_inside.chocolate.led <= red;
    machine_info_inside.chocolate.monitor <= 10'd0;
    machine_info_inside.froth.led <= red;
    machine_info_inside.froth.monitor <= 10'd0;
    machine_flavor_out = no_coffee;

    #5;
    inf.rst_n  <= 1;
    $display("*************************");
    $display("**** Finish RESET    ****");
    $display("*************************");
end
endtask

//------------------Input Supply----------------------
task input_supply(logic full);
begin
    machine_flavor_out = no_coffee;
    if (full == 0) begin
        repeat(1) @(negedge clk);
        i = supply_input_rand.randomize();
        
        supply_limit = 1023 - machine_info_inside.espresso.monitor;
        if (supply_input_rand.espresso == 1'd1) begin
            if (supply_limit >= supply_input_rand.e_supply_amount) begin
                inf.select_i <= espresso;
                inf.supply <= supply_input_rand.e_supply_amount;
                machine_info_inside.espresso.monitor += supply_input_rand.e_supply_amount;
                repeat(1) @(negedge clk);
            end else begin 
                if (supply_limit !== 0) begin
                    inf.select_i <= espresso;
                    inf.supply <= supply_limit;
                    machine_info_inside.espresso.monitor += supply_limit;
                    repeat(1) @(negedge clk);
                end
            end
        end

        supply_limit = 1023 - machine_info_inside.milk.monitor;
        if (supply_input_rand.milk == 1'd1) begin
            if (supply_limit >= supply_input_rand.m_supply_amount) begin
                inf.select_i <= milk;
                inf.supply <= supply_input_rand.m_supply_amount;
                machine_info_inside.milk.monitor += supply_input_rand.m_supply_amount;
                repeat(1) @(negedge clk);
            end else begin 
                if (supply_limit !== 0) begin
                    inf.select_i <= milk;
                    inf.supply <= supply_limit;
                    machine_info_inside.milk.monitor += supply_limit;
                    repeat(1) @(negedge clk);
                end
            end
        end

        supply_limit = 1023 - machine_info_inside.chocolate.monitor;
        if (supply_input_rand.chocolate == 1'd1) begin
            if (supply_limit >= supply_input_rand.c_supply_amount) begin
                inf.select_i <= chocolate;
                inf.supply <= supply_input_rand.c_supply_amount;
                machine_info_inside.chocolate.monitor += supply_input_rand.c_supply_amount;
                repeat(1) @(negedge clk);
            end else begin 
                if (supply_limit !== 0) begin
                    inf.select_i <= chocolate;
                    inf.supply <= supply_limit;
                    machine_info_inside.chocolate.monitor += supply_limit;
                    repeat(1) @(negedge clk);
                end
            end
        end

        supply_limit = 1023 - machine_info_inside.froth.monitor;
        if (supply_input_rand.froth == 1'd1) begin
            if (supply_limit >= supply_input_rand.f_supply_amount) begin
                inf.select_i <= froth;
                inf.supply <= supply_input_rand.f_supply_amount;
                machine_info_inside.froth.monitor += supply_input_rand.f_supply_amount;
                repeat(1) @(negedge clk);
            end else begin 
                if (supply_limit !== 0) begin
                    inf.select_i <= froth;
                    inf.supply <= supply_limit;
                    machine_info_inside.froth.monitor += supply_limit;
                    repeat(1) @(negedge clk);
                end
            end
        end
    end else begin
        repeat(1) @(negedge clk);
        i = supply_input_rand.randomize();
        
        supply_limit = 1023 - machine_info_inside.espresso.monitor;
        if (supply_limit !== 0) begin
            inf.select_i <= espresso;
            inf.supply <= supply_limit;
            machine_info_inside.espresso.monitor += supply_limit;
            repeat(1) @(negedge clk);
        end
        supply_limit = 1023 - machine_info_inside.milk.monitor;
        if (supply_limit !== 0) begin
            inf.select_i <= milk;
            inf.supply <= supply_limit;
            machine_info_inside.milk.monitor += supply_limit;
            repeat(1) @(negedge clk);
        end
        supply_limit = 1023 - machine_info_inside.chocolate.monitor;
        if (supply_limit !== 0) begin
            inf.select_i <= chocolate;
            inf.supply <= supply_limit;
            machine_info_inside.chocolate.monitor += supply_limit;
            repeat(1) @(negedge clk);
        end
        supply_limit = 1023 - machine_info_inside.froth.monitor;
        if (supply_limit !== 0) begin
            inf.select_i <= froth;
            inf.supply <= supply_limit;
            machine_info_inside.froth.monitor += supply_limit;
            repeat(1) @(negedge clk);
        end
    end

    if (machine_info_inside.espresso.monitor > 0) 
        machine_info_inside.espresso.led = green;
    else 
        machine_info_inside.espresso.led = red;

    if (machine_info_inside.milk.monitor > 0) 
        machine_info_inside.milk.led = green;
    else 
        machine_info_inside.milk.led = red;

    if (machine_info_inside.chocolate.monitor > 0) 
        machine_info_inside.chocolate.led = green;
    else 
        machine_info_inside.chocolate.led = red;

    if (machine_info_inside.froth.monitor > 0) 
        machine_info_inside.froth.led = green;
    else 
        machine_info_inside.froth.led = red;

    inf.select_i <= none;
    inf.supply <= 10'd0;
    repeat(1)@(negedge clk);

    out_valid_check();
    window_check();
    flavor_out_check();
    out_valid_one_cycle();
end
endtask

//-----------Press Button & Check-------------
task press_buttom(select_flavor select_flavor_rand,
                  select_size select_size_rand,
                  select_ratio select_ratio_rand);
begin

    if (select_flavor_rand.flavor_in == user_define) begin
        inf.flavor_btn <= select_flavor_rand.flavor_in;
        inf.required_size <= select_size_rand.size_in;
        inf.ratio <= select_ratio_rand.espresso;
        repeat(1)@(negedge clk);

        inf.flavor_btn <= no_coffee;
        inf.required_size <= no_size_inf;
        inf.ratio <= select_ratio_rand.milk;
        repeat(1)@(negedge clk);

        inf.ratio <= select_ratio_rand.chocolate;
        repeat(1)@(negedge clk);

        inf.ratio <= select_ratio_rand.froth;
        repeat(1)@(negedge clk);

    end else begin
        inf.flavor_btn <= select_flavor_rand.flavor_in;
        inf.required_size <= select_size_rand.size_in;
        repeat(1)@(negedge clk);

    end

    // calculate solution
    gcd = 1;
    for (i = 2; i < 8; i++) begin
        if (select_ratio_rand.espresso % i == 0 &&
            select_ratio_rand.milk % i == 0 &&
            select_ratio_rand.chocolate % i == 0 &&
            select_ratio_rand.froth % i == 0)
            gcd = i; 
    end

    case (select_size_rand.size_in)
        s: capacity = 240;
        m: capacity = 360;
        l: capacity = 480;
        xl: capacity = 600;
        default: capacity = 0;
    endcase

    total_ratio = (select_ratio_rand.espresso +
                   select_ratio_rand.milk + 
                   select_ratio_rand.chocolate +
                   select_ratio_rand.froth) / gcd; 

    case (select_flavor_rand.flavor_in)
        latte: 
            begin
                required_espresso = capacity / 10 * 3;
                required_milk = capacity / 10 * 3;
                required_chocolate = 0;
                required_froth = capacity / 10 * 4;
            end
        cappuccino: 
            begin
                required_espresso = capacity / 15 * 7;
                required_milk = capacity / 15 * 3;
                required_chocolate = 0;
                required_froth = capacity / 15 * 5;
            end
        mocha: 
            begin
                required_espresso = capacity / 5 * 3;
                required_milk = capacity / 5;
                required_chocolate = capacity / 5 ;
                required_froth = 0;
            end
        user_define:
            begin
                required_espresso = capacity / total_ratio * (select_ratio_rand.espresso / gcd);
                required_milk = capacity / total_ratio * (select_ratio_rand.milk / gcd);
                required_chocolate = capacity / total_ratio * (select_ratio_rand.chocolate / gcd); 
                required_froth = capacity / total_ratio * (select_ratio_rand.froth / gcd);
            end
        default:
            begin
                required_espresso = 0;
                required_milk = 0;
                required_chocolate = 0;
                required_froth = 0;
            end
    endcase

    if (machine_info_inside.espresso.monitor >= required_espresso &&
        machine_info_inside.milk.monitor >= required_milk &&
        machine_info_inside.chocolate.monitor >= required_chocolate &&
        machine_info_inside.froth.monitor >= required_froth) begin

        machine_info_inside.espresso.monitor -= required_espresso;
        machine_info_inside.milk.monitor -= required_milk;
        machine_info_inside.chocolate.monitor -= required_chocolate;
        machine_info_inside.froth.monitor -= required_froth;
        machine_flavor_out = select_flavor_rand.flavor_in;

        if (machine_info_inside.espresso.monitor > 0) 
            machine_info_inside.espresso.led = green;
        else 
            machine_info_inside.espresso.led = red;

        if (machine_info_inside.milk.monitor > 0) 
            machine_info_inside.milk.led = green;
        else 
            machine_info_inside.milk.led = red;

        if (machine_info_inside.chocolate.monitor > 0) 
            machine_info_inside.chocolate.led = green;
        else 
            machine_info_inside.chocolate.led = red;

        if (machine_info_inside.froth.monitor > 0) 
            machine_info_inside.froth.led = green;
        else 
            machine_info_inside.froth.led = red;

    end else begin
        machine_flavor_out = no_coffee;
        if (required_espresso > machine_info_inside.espresso.monitor ||
            machine_info_inside.espresso.monitor == 0)
            machine_info_inside.espresso.led = red;
        else
            machine_info_inside.espresso.led = green;

        if (required_milk > machine_info_inside.milk.monitor ||
            machine_info_inside.milk.monitor == 0)
            machine_info_inside.milk.led = red;
        else
            machine_info_inside.milk.led = green;

        if (required_chocolate > machine_info_inside.chocolate.monitor ||
            machine_info_inside.chocolate.monitor == 0)
            machine_info_inside.chocolate.led = red;
        else
            machine_info_inside.chocolate.led = green;

        if (required_froth > machine_info_inside.froth.monitor ||
            machine_info_inside.froth.monitor == 0)
            machine_info_inside.froth.led = red;
        else
            machine_info_inside.froth.led = green;
    end


    inf.ratio <= 3'd0;
    inf.flavor_btn <= no_coffee;
    inf.required_size <= no_size_inf;
    repeat(1)@(negedge clk);

    out_valid_check();
    window_check();
    flavor_out_check();
    out_valid_one_cycle();

    // after press button
    machine_flavor_out = no_coffee;
end
endtask

//-----------Checkt out_valid---------------
task out_valid_check(); begin
    check_output_times = 0;
    while(inf.out_valid !== 1 && check_output_times < 30) begin
	check_output_times = check_output_times + 1;
	repeat(1)@(negedge clk);
    end
    if(check_output_times == 30) begin
	$display("-----Your out_valid should be high in 30 cycles------\n");
        fail;
    end
end
endtask

task out_valid_one_cycle(); begin
    repeat(1)@(negedge clk);
    if(inf.out_valid) begin
        $display("-----Your out_valid should be high onlu one cycle------\n");
        fail;
    end
end
endtask

//-----------Check window value-----------------
task window_check();
begin
    if((inf.window.espresso.led !== machine_info_inside.espresso.led) ||
       (inf.window.espresso.monitor !== machine_info_inside.espresso.monitor)) begin
            $display("-------Espresso Window Wrong------- at time: %t",$time);
            $display("Gold led:%d, Your led: %d",
                machine_info_inside.espresso.led,
                inf.window.espresso.led);
            $display("Gold Monitor:%d, Your Monitor: %d",
                machine_info_inside.espresso.monitor,
                inf.window.espresso.monitor);
            fail;
    end

    if((inf.window.milk.led !== machine_info_inside.milk.led) ||
       (inf.window.milk.monitor !== machine_info_inside.milk.monitor)) begin
            $display("-------Milk Window Wrong------- at time: %t",$time);
            $display("Gold led:%d, Your led: %d",
                machine_info_inside.milk.led,
                inf.window.milk.led);
            $display("Gold Monitor:%d, Your Monitor: %d",
                machine_info_inside.milk.monitor,
                inf.window.milk.monitor);
            fail;
    end

    if((inf.window.chocolate.led !== machine_info_inside.chocolate.led) ||
       (inf.window.chocolate.monitor !== machine_info_inside.chocolate.monitor)) begin
            $display("-------Chocolate Window Wrong------- at time: %t",$time);
            $display("Gold led:%d, Your led: %d",
                machine_info_inside.chocolate.led,
                inf.window.chocolate.led);
            $display("Gold Monitor:%d, Your Monitor: %d",
                machine_info_inside.chocolate.monitor,
                inf.window.chocolate.monitor);
            fail;
    end

    if((inf.window.froth.led !== machine_info_inside.froth.led) ||
       (inf.window.froth.monitor !== machine_info_inside.froth.monitor)) begin
            $display("-------Froth Window Wrong------- at time: %t",$time);
            $display("Gold led:%d, Your led: %d",
                machine_info_inside.froth.led,
                inf.window.froth.led);
            $display("Gold Monitor:%d, Your Monitor: %d",
                machine_info_inside.froth.monitor,
                inf.window.froth.monitor);
            fail;
    end
end
endtask

//-----------Check flavor_out----------------
task flavor_out_check;
begin
    if(inf.flavor_out !== machine_flavor_out) begin
        $display("-------flavor_out Wrong-------%t",$time);
        $display("Gold flavor_out: %d , not %d",
            machine_flavor_out,
            inf.flavor_out);
	fail;
    end	
end
endtask


task fail;
begin
	repeat(10)@(negedge clk);

	$display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOoooooo888888OOOOOOOOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOO88OOoc:.                   cOOOOOOOOOOOOOOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOOOOOOOOOO8O.                             oOOOOOOOOOOOOOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOOOOOO8O.                                     oOOOOOOOOOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOOOOO:                                            O8OOOOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOO8c                                                 O8OOOOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOO8.                                                     O8OOOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOO8.                                                         8OOOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOc                                                            oOOOOOOOOOOOOO");
	$display("OOOOOOOOOO8c                                                              C8OOOOOOOOOOO");
	$display("OOOOOOOOO8                                                                 .OOOOOOOOOOO");
	$display("OOOOOOOOO.                                                                  c8OOOOOOOOO");
	$display("OOOOOOO8                                                                      8OOOOOOOO");
	$display("OOOOOOO:                      C.            :.            O@                  o8OOOOOOO");
	$display("OOOOO8.                      O@@C          o@@8:        C@@@@C                 oOOOOOOO");
	$display("OOOOOO          :O         .@@@@@@o       @@@@@@@C    8@@@@@@@8.        8:      8OOOOOO");
	$display("OOOOO          .@@@@      @@@@@@@@@@C   @@@@@@@@@@@@@@@@@@@@@@@@O.    @@@@o     o8OOOOO");
	$display("OOOO.         C@@@@@@@:.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:C@@@@@@@@@@@@@@@@@@@@.    COOOOO");
	$display("OOO8    .@    @@@@@@@@@@@@@@O@@@@@@@@@@@@@@@@@@@@@@@@@  .O@@@@@@@@@@@@@@@@@@@O    OOOOO");
	$display("OO8O    @@@@@@@@@@@@@@@@@@  @@@@@@@@@@@@@@@@@@@@@@@@@@@o       .:cCo  @@@@@@@@C   OOOOO");
	$display("OO8o   C@@@@@@@@@@@@@@@c  :@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@O8OOoCO@@@@@@@@@@@@@@  c8OOO");
	$display("OOO:  C@@@@@@c          c@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@8.       cO@@@@@@@@@@@@  .OOOO");
	$display("OOO.  @@@@@@@@@8c:coC8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:   OO          :8@@@@@@@@.  oOOO");
	$display("OOO   @@@@@@@@@8.           .o@@@@@@o c@@@@@@@@@@@@@: .O@@@C      @@@O  .8@@@@@@.  oOOO");
	$display("OOO   @@@@@@@o   cO       @O:   8@@@@: c@@@@@@@@@@@@                      8@@@@@.  oOOO");
	$display("OOO.  @@@@@@  c@@@@c      .     .8@@C:  @@@@@@@@@@@@@@8OoooCOO8@@@@8OOooO@@@@@@@.  oOOO");
	$display("OOO.  8@@@@:              coOO@@@8    co@@@@@@@@@@@@@@@@@@@@@@@8      ..@@@@@@@@.  oOOO");
	$display("OOO:  o@@@@@@@@@@@@@@@8C8@@@@@@@@@   :@@@@@@@@@@@@@@@@...... .@@@@@@@@OC@@@@@@@@.  oOOO");
	$display("OO8O   O@@@@@@@@8       C@@@@@@@@@@@   O@@@@@@@@@@@@@@Cooo    C@@@@@@@@@@@@@@@@@   COOO");
	$display("OOO8   o@@@@@@@@8::cO8@@@@@@@@@@@@@@@O8@@@@@@@@@@@@@@@@@O     .8@@@@@@@@@@@@@@@@   OOOO");
	$display("OOO8.   @@@@@@@@@@@@@@@@Oo    @@@@@@@@@@@@@@@@@@@@@@@@@c  C@C  .@@@@@@@@@@@@@@@@  c8OOO");
	$display("OOOOC   8@@@@@@@@@@@@@8    o@@@@@@@@@@@@@@@@@@@@@@@@@C  .@@@@8  @@@@@@@@@@@@@@@:  O8OOO");
	$display("OOOO8o  .@@@@@@@@@@@@@@O  .   o@@@@@@@@@@@@@@@@@@@8c   O@@@@@@@@@@@@@@@@@@@@@@:   8OOOO");
	$display("OOOOO8   .@@@@@@@@@@@@@@  O@8o    :o8@@@@@@@@@Oo    .8@@@@@@@@@@@@@@@@@@@@@@@@   oOOOOO");
	$display("OOOOOOc   8@@@@@@@@@@@@@@@@@@@@@Oo                 o@@@@@@@@@@@@@@@@@@@@@@@@8.  o8OOOOO");
	$display("OOOOOO8o   o@@@@@@@@@@@@@@@@@@@@@@@@c   C@@@@@:  c@@@@@@@@@@@@@@@@@@@@@@@@@@    8OOOOOO");
	$display("OOOOOOO8    @@@@@@@@@@@@@@@@@@@@@@@@@@@@.     .O@@@@@@@@@@@@@@@@@@@@@@@@@@@:  c8OOOOOOO");
	$display("OOOOOOOOOc   8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@C. .@@@@@@@@@@@@@@@@@@@@@@@@    8OOOOOOOO");
	$display("OOOOOOOOO8.   @@@@@@@@@@@@@@@@@@@@@@@@@@@@     .@@@@@@@@@@@@@@@@@@@@@@@@.   c8OOOOOOOOO");
	$display("OOOOOOOOOO8C   .@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@o    COOOOOOOOOOO");
	$display("OOOOOOOOOOOOC    o@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@o   .COOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOO.   c@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:      COOOOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOo    8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@O    O@8c  C8OOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOOOC.      O@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@8C     c@C  @8:   OOOOOOOOOOO");
	$display("OOOOOOOOOOOOOOOOO8  .8         .oO@@@@@@@@@@@@@@@@@@8O:      c888888o  C8O  :8OOOOOOOOO");
	$display("OOOOOOOOOOOOOOOO8c  88 .  ....                          oO888888888888  88c   8OOOOOOOO");
	$display("OOOOOOOOOOOOOOOO.   @:.8.   ....  C@@8OOoocccoooO888888888888888888888O  C@C  8OOOOOOOO");

	$display("fail");
	$finish;
end
endtask

task pass;
begin
	$display("\n");
	$display("88888888888888888888888                             888888888888888888888");
	$display("8888888888888888888888                                8C88888888888888888");
	$display("88888888888888888C.                                    o88888888888888888");
	$display("888888888888888C.                                         C88888888888888");
	$display("888888888888                                                C888888888888");
	$display("8888888888o                                                  .O8888888888");
	$display("88888888O                                                      :888888888");
	$display("8888888                                                          O8888888");
	$display("888888c                                                           o888888");
	$display("88888:           @C                 c:                             o88888");
	$display("888O. o      :8@@@@@@O           @@@@@@:          c@@@@8.           :8888");
	$display("888: c@     @@@@@@@@@@@.      o@@@@@@@@@@c     :@@@@@@@@@O      .o:  8888");
	$display("88. c@@@Oc.    .c@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:.C@@@@@C c888");
	$display("88  @@o c8@@@@@@8  o@@@@@@@@@@@@@@@@@@@@@@@@@@C:      O@@@@@@@@@@@@@. O88");
	$display("88 cO :@@@@@@@@@@@@. C@@@@@@@@@@@@@@@@@@@@@.  o8@@@@@@c  c@@@@@@@@@@o c88");
	$display("8O  c@@@C       :@@@@: @@@@@@@@@@@@@@@@@@c @@@@@@@@@@@@@@8 C@@@@@@@@8  O8");
	$display("8C .@@@.         :@@@@ @@@@@@@@@@@@@@@@@. 8@@@o       @@@@@ c@@@@@@@@  C8");
	$display("8o C@@@   c@@@c   o@@@cC@@@@@@@@@@@@@@@  @@@c           8@@o o@@@@@@@  o8");
	$display("8C o@@@   :@@@.   O@@@:O@@@@@@@@@@@@@@O c@@8    @@@8    c@@O :@@@@@@@  c8");
	$display("8C  @@@c         c@@@C @@@@@@@@@@@@@@@O :@@8    @@@@:   o@@O :@@@@@@@  C8");
	$display("8O   :@@@@8o.:o8@@@O  O@@O 8@@@@@@@@@@@: C@@8          c@@@  @@@@@@@O .88");
	$display("C8 :O  C@@@@@@@@@o  o@@    @@@@@@@@@@@@@  o@@@O:      @@@@O 8@@@@@@@c C88");
	$display("88  O@@:    .    :8@@@@ 8@@@@@@@@@@@@@@@@: O@@@@@@@@@@@@8. @@@@@@@@8 :888");
	$display("OC   o@@@@@@@@@@@@8:O@@@8@@@@@@@@@: O@@@@@@O:   ::::   .C@@@@@@@@@8  8C88");
	$display("@8o   o@@@@@@@@@@@ :@@@@@@@@@8Oo:     @@@@@@@@@@8888@@@@@@@@@@@@@8     O@");
	$display("@@8OO. O@@@@@@@@@@@@.:@@  8@@  C@c  :@@@@@@@@@@@@@@@@@@@@@@@@@@@o    @@@@");
	$display("@@@@OOc c@@@@@@@@@@@O \033[91m  c. : .C:.c. \033[0mO@@@@@@@@@@@@@@@@@@@@@@@@@@@   C@@@@O");
	$display("C@@@@8O  .@@@@@@@@@@@@@\033[91m oOOOOOOOOC \033[0m:@@@@@@@@@@@@@@@@@@@@@@@@@@@. o@@@@8OO");
	$display("08@@@@@    .@@@@@@@@@@@@.\033[91m COOOOOO \033[0m.@@@@@@@@@@@@@@@@@@@@@@@@@:  . C@@8OO88");
	$display("888@@@oo@8. .8@@@@@@@@@@@:\033[91m COOOOO \033[0m@@@@@@@@@@@@@@@@@@@@@@@@o  .O8O0:COC00O");
	$display("880co0o88888:   o@@@@@@@@@@\033[91m COOC \033[0m@@@@@@@@@@@@@@@@@@@@@c   .@88888@o088O88");
	$display("88C0888888888Oc   .O@@@@@@@@\033[91m :O. \033[0m@@@@@@@@@@@@@@@@@@8c   c888888CC@8O08888");
	$display("8808888888CO888OCc.   c@@@@@@.  O@@@@@@@@@@@@@@@:     O88888888800O@80O88");
	$display("O0O8888888888c8888OCCCC     cCOO8@8OOOCoc:.     cCO88888888888CC8@888888O");
	$display("8888888C@OC8888888888OCCCCoc.             .coCCO88888888888888cCCC8888880");
	$display("-------------------------------------------");
	$display("Awesome!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!");
	$display("You Pass Lab09!!!!!!!!!!!!!!!!!!!!!!!!!!!!!");
	$display("-------------------------------------------");
	$timeformat(-9, 5, " ns", 10); 
        $display("Your total simulation time = %t", $time);
	$write("\033[0m ");
	$finish;
end
endtask
endprogram
